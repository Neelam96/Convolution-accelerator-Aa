-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accMemAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    acc_mem_request_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    acc_mem_request_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    acc_mem_request_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    acc_mem_response_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    acc_mem_response_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    acc_mem_response_1_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accMemAccessDaemon;
architecture accMemAccessDaemon_arch of accMemAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal accMemAccessDaemon_CP_248_start: Boolean;
  signal accMemAccessDaemon_CP_248_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_82_branch_req_0 : boolean;
  signal RPIPE_acc_mem_request_1_85_inst_req_0 : boolean;
  signal RPIPE_acc_mem_request_1_85_inst_ack_0 : boolean;
  signal RPIPE_acc_mem_request_1_85_inst_req_1 : boolean;
  signal RPIPE_acc_mem_request_1_85_inst_ack_1 : boolean;
  signal call_stmt_108_call_req_0 : boolean;
  signal call_stmt_108_call_ack_0 : boolean;
  signal call_stmt_108_call_req_1 : boolean;
  signal call_stmt_108_call_ack_1 : boolean;
  signal WPIPE_acc_mem_response_1_109_inst_req_0 : boolean;
  signal WPIPE_acc_mem_response_1_109_inst_ack_0 : boolean;
  signal WPIPE_acc_mem_response_1_109_inst_req_1 : boolean;
  signal WPIPE_acc_mem_response_1_109_inst_ack_1 : boolean;
  signal do_while_stmt_82_branch_ack_0 : boolean;
  signal do_while_stmt_82_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accMemAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accMemAccessDaemon_CP_248_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accMemAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_248_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_248_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accMemAccessDaemon_CP_248_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accMemAccessDaemon_CP_248_start,"accMemAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accMemAccessDaemon_CP_248_symbol, "accMemAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accMemAccessDaemon_CP_248: Block -- control-path 
    signal accMemAccessDaemon_CP_248_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    accMemAccessDaemon_CP_248_elements(0) <= accMemAccessDaemon_CP_248_start;
    accMemAccessDaemon_CP_248_symbol <= accMemAccessDaemon_CP_248_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_81/$entry
      -- CP-element group 0: 	 branch_block_stmt_81/branch_block_stmt_81__entry__
      -- CP-element group 0: 	 branch_block_stmt_81/do_while_stmt_82__entry__
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	24 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_81/$exit
      -- CP-element group 1: 	 branch_block_stmt_81/branch_block_stmt_81__exit__
      -- CP-element group 1: 	 branch_block_stmt_81/do_while_stmt_82__exit__
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(1) <= accMemAccessDaemon_CP_248_elements(24);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_81/do_while_stmt_82/$entry
      -- CP-element group 2: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82__entry__
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(2) <= accMemAccessDaemon_CP_248_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	24 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82__exit__
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accMemAccessDaemon_CP_248_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_81/do_while_stmt_82/loop_back
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accMemAccessDaemon_CP_248_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: 	23 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_81/do_while_stmt_82/condition_done
      -- CP-element group 5: 	 branch_block_stmt_81/do_while_stmt_82/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_81/do_while_stmt_82/loop_taken/$entry
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(5) <= accMemAccessDaemon_CP_248_elements(21);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	20 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_81/do_while_stmt_82/loop_body_done
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(6) <= accMemAccessDaemon_CP_248_elements(20);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(7) <= accMemAccessDaemon_CP_248_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(8) <= accMemAccessDaemon_CP_248_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/loop_body_start
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accMemAccessDaemon_CP_248_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Sample/rr
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:RPIPE_acc_mem_request_1_85_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(10), ack => RPIPE_acc_mem_request_1_85_inst_req_0); -- 
    accMemAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accMemAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accMemAccessDaemon_CP_248_elements(9) & accMemAccessDaemon_CP_248_elements(13);
      gj_accMemAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_update_start_
      -- CP-element group 11: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Update/cr
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:RPIPE_acc_mem_request_1_85_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(11), ack => RPIPE_acc_mem_request_1_85_inst_req_1); -- 
    accMemAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accMemAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accMemAccessDaemon_CP_248_elements(12) & accMemAccessDaemon_CP_248_elements(16);
      gj_accMemAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Sample/ra
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:RPIPE_acc_mem_request_1_85_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_acc_mem_request_1_85_inst_ack_0, ack => accMemAccessDaemon_CP_248_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/RPIPE_acc_mem_request_1_85_Update/ca
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:RPIPE_acc_mem_request_1_85_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_acc_mem_request_1_85_inst_ack_1, ack => accMemAccessDaemon_CP_248_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Sample/crr
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_108_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(14), ack => call_stmt_108_call_req_0); -- 
    accMemAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accMemAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accMemAccessDaemon_CP_248_elements(13) & accMemAccessDaemon_CP_248_elements(16);
      gj_accMemAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_update_start_
      -- CP-element group 15: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Update/ccr
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_108_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(15), ack => call_stmt_108_call_req_1); -- 
    accMemAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "accMemAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accMemAccessDaemon_CP_248_elements(19);
      gj_accMemAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Sample/cra
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_108_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_108_call_ack_0, ack => accMemAccessDaemon_CP_248_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/call_stmt_108_Update/cca
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:call_stmt_108_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_108_call_ack_1, ack => accMemAccessDaemon_CP_248_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Sample/req
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:WPIPE_acc_mem_response_1_109_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(18), ack => WPIPE_acc_mem_response_1_109_inst_req_0); -- 
    accMemAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accMemAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accMemAccessDaemon_CP_248_elements(17) & accMemAccessDaemon_CP_248_elements(20);
      gj_accMemAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_update_start_
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Update/req
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:WPIPE_acc_mem_response_1_109_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:WPIPE_acc_mem_response_1_109_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_response_1_109_inst_ack_0, ack => accMemAccessDaemon_CP_248_elements(19)); -- 
    req_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(19), ack => WPIPE_acc_mem_response_1_109_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (4) 
      -- CP-element group 20: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/$exit
      -- CP-element group 20: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/WPIPE_acc_mem_response_1_109_Update/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:WPIPE_acc_mem_response_1_109_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_acc_mem_response_1_109_inst_ack_1, ack => accMemAccessDaemon_CP_248_elements(20)); -- 
    -- CP-element group 21:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	5 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/condition_evaluated
      -- CP-element group 21: 	 branch_block_stmt_81/do_while_stmt_82/do_while_stmt_82_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:do_while_stmt_82_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accMemAccessDaemon_CP_248_elements(21), ack => do_while_stmt_82_branch_req_0); -- 
    -- Element group accMemAccessDaemon_CP_248_elements(21) is a control-delay.
    cp_element_21_delay: control_delay_element  generic map(name => " 21_delay", delay_value => 1)  port map(req => accMemAccessDaemon_CP_248_elements(9), ack => accMemAccessDaemon_CP_248_elements(21), clk => clk, reset =>reset);
    -- CP-element group 22:  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_81/do_while_stmt_82/loop_exit/$exit
      -- CP-element group 22: 	 branch_block_stmt_81/do_while_stmt_82/loop_exit/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:do_while_stmt_82_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_82_branch_ack_0, ack => accMemAccessDaemon_CP_248_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	5 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_81/do_while_stmt_82/loop_taken/$exit
      -- CP-element group 23: 	 branch_block_stmt_81/do_while_stmt_82/loop_taken/ack
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:do_while_stmt_82_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_82_branch_ack_1, ack => accMemAccessDaemon_CP_248_elements(23)); -- 
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	3 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	1 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_81/do_while_stmt_82/$exit
      -- 
    -- logger for CP element group accMemAccessDaemon_CP_248_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accMemAccessDaemon_CP_248_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accMemAccessDaemon:CP:accMemAccessDaemon_CP_248_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    accMemAccessDaemon_CP_248_elements(24) <= accMemAccessDaemon_CP_248_elements(3);
    accMemAccessDaemon_do_while_stmt_82_terminator_325: loop_terminator -- 
      generic map (name => " accMemAccessDaemon_do_while_stmt_82_terminator_325", max_iterations_in_flight =>20) 
      port map(loop_body_exit => accMemAccessDaemon_CP_248_elements(6),loop_continue => accMemAccessDaemon_CP_248_elements(23),loop_terminate => accMemAccessDaemon_CP_248_elements(22),loop_back => accMemAccessDaemon_CP_248_elements(4),loop_exit => accMemAccessDaemon_CP_248_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_273_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= accMemAccessDaemon_CP_248_elements(7);
        preds(1)  <= accMemAccessDaemon_CP_248_elements(8);
        entry_tmerge_273 : transition_merge -- 
          generic map(name => " entry_tmerge_273")
          port map (preds => preds, symbol_out => accMemAccessDaemon_CP_248_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal cmd_1_86 : std_logic_vector(31 downto 0);
    signal col_index1_98 : std_logic_vector(4 downto 0);
    signal konst_113_wire_constant : std_logic_vector(0 downto 0);
    signal rdata1_108 : std_logic_vector(15 downto 0);
    signal row_index1_94 : std_logic_vector(5 downto 0);
    signal rwbar1_102 : std_logic_vector(0 downto 0);
    signal wdata1_90 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    konst_113_wire_constant <= "1";
    -- logger for split-operator slice_101_inst flow-through 
    process(rwbar1_102) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_101_inst:flowthrough inputs: " & " cmd_1_86 = "& Convert_SLV_To_Hex_String(cmd_1_86) & " outputs:" & " rwbar1_102= "  & Convert_SLV_To_Hex_String(rwbar1_102));
      --
    end process; 
    -- flow-through slice operator slice_101_inst
    rwbar1_102 <= cmd_1_86(0 downto 0);
    -- logger for split-operator slice_89_inst flow-through 
    process(wdata1_90) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_89_inst:flowthrough inputs: " & " cmd_1_86 = "& Convert_SLV_To_Hex_String(cmd_1_86) & " outputs:" & " wdata1_90= "  & Convert_SLV_To_Hex_String(wdata1_90));
      --
    end process; 
    -- flow-through slice operator slice_89_inst
    wdata1_90 <= cmd_1_86(31 downto 16);
    -- logger for split-operator slice_93_inst flow-through 
    process(row_index1_94) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_93_inst:flowthrough inputs: " & " cmd_1_86 = "& Convert_SLV_To_Hex_String(cmd_1_86) & " outputs:" & " row_index1_94= "  & Convert_SLV_To_Hex_String(row_index1_94));
      --
    end process; 
    -- flow-through slice operator slice_93_inst
    row_index1_94 <= cmd_1_86(15 downto 10);
    -- logger for split-operator slice_97_inst flow-through 
    process(col_index1_98) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:slice_97_inst:flowthrough inputs: " & " cmd_1_86 = "& Convert_SLV_To_Hex_String(cmd_1_86) & " outputs:" & " col_index1_98= "  & Convert_SLV_To_Hex_String(col_index1_98));
      --
    end process; 
    -- flow-through slice operator slice_97_inst
    col_index1_98 <= cmd_1_86(9 downto 5);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_82_branch_req_0," req0 do_while_stmt_82_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_82_branch_ack_0," ack0 do_while_stmt_82_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_82_branch_ack_1," ack1 do_while_stmt_82_branch");
    do_while_stmt_82_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_113_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_82_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_82_branch_req_0,
          ack0 => do_while_stmt_82_branch_ack_0,
          ack1 => do_while_stmt_82_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_acc_mem_request_1_85_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_acc_mem_request_1_85_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:RPIPE_acc_mem_request_1_85_inst:started:   PipeRead from acc_mem_request_1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_acc_mem_request_1_85_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:RPIPE_acc_mem_request_1_85_inst:finished:  outputs: " & " cmd_1_86= "  & Convert_SLV_To_Hex_String(cmd_1_86));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_acc_mem_request_1_85_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_acc_mem_request_1_85_inst_req_0;
      RPIPE_acc_mem_request_1_85_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_acc_mem_request_1_85_inst_req_1;
      RPIPE_acc_mem_request_1_85_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_1_86 <= data_out(31 downto 0);
      acc_mem_request_1_read_0_gI: SplitGuardInterface generic map(name => "acc_mem_request_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      acc_mem_request_1_read_0: InputPortRevised -- 
        generic map ( name => "acc_mem_request_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => acc_mem_request_1_pipe_read_req(0),
          oack => acc_mem_request_1_pipe_read_ack(0),
          odata => acc_mem_request_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_acc_mem_response_1_109_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_acc_mem_response_1_109_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:WPIPE_acc_mem_response_1_109_inst:started:   PipeWrite to acc_mem_response_1 inputs: " & " rdata1_108 = "& Convert_SLV_To_Hex_String(rdata1_108));
          --
        end if; 
        if WPIPE_acc_mem_response_1_109_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:WPIPE_acc_mem_response_1_109_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_acc_mem_response_1_109_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_acc_mem_response_1_109_inst_req_0;
      WPIPE_acc_mem_response_1_109_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_acc_mem_response_1_109_inst_req_1;
      WPIPE_acc_mem_response_1_109_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata1_108;
      acc_mem_response_1_write_0_gI: SplitGuardInterface generic map(name => "acc_mem_response_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      acc_mem_response_1_write_0: OutputPortRevised -- 
        generic map ( name => "acc_mem_response_1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => acc_mem_response_1_pipe_write_req(0),
          oack => acc_mem_response_1_pipe_write_ack(0),
          odata => acc_mem_response_1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_108_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_108_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:call_stmt_108_call:started:  Call to module accessMem inputs: " & " rwbar1_102 = "& Convert_SLV_To_Hex_String(rwbar1_102) & " row_index1_94 = "& Convert_SLV_To_Hex_String(row_index1_94) & " col_index1_98 = "& Convert_SLV_To_Hex_String(col_index1_98) & " wdata1_90 = "& Convert_SLV_To_Hex_String(wdata1_90));
          --
        end if; 
        if call_stmt_108_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accMemAccessDaemon:DP:call_stmt_108_call:finished:  outputs: " & " rdata1_108= "  & Convert_SLV_To_Hex_String(rdata1_108));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_108_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_108_call_req_0;
      call_stmt_108_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_108_call_req_1;
      call_stmt_108_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar1_102 & row_index1_94 & col_index1_98 & wdata1_90;
      rdata1_108 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 28,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 5,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end accMemAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accelerator is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_accelerator_pipe_read_req : out  std_logic_vector(0 downto 0);
    start_accelerator_pipe_read_ack : in   std_logic_vector(0 downto 0);
    start_accelerator_pipe_read_data : in   std_logic_vector(15 downto 0);
    accelerator_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    accelerator_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    accelerator_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    read_sums_pipe_write_req : out  std_logic_vector(0 downto 0);
    read_sums_pipe_write_ack : in   std_logic_vector(0 downto 0);
    read_sums_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    initIfMaps_call_reqs : out  std_logic_vector(0 downto 0);
    initIfMaps_call_acks : in   std_logic_vector(0 downto 0);
    initIfMaps_call_data : out  std_logic_vector(13 downto 0);
    initIfMaps_call_tag  :  out  std_logic_vector(0 downto 0);
    initIfMaps_return_reqs : out  std_logic_vector(0 downto 0);
    initIfMaps_return_acks : in   std_logic_vector(0 downto 0);
    initIfMaps_return_data : in   std_logic_vector(1 downto 0);
    initIfMaps_return_tag :  in   std_logic_vector(0 downto 0);
    initFilter_call_reqs : out  std_logic_vector(0 downto 0);
    initFilter_call_acks : in   std_logic_vector(0 downto 0);
    initFilter_call_data : out  std_logic_vector(5 downto 0);
    initFilter_call_tag  :  out  std_logic_vector(0 downto 0);
    initFilter_return_reqs : out  std_logic_vector(0 downto 0);
    initFilter_return_acks : in   std_logic_vector(0 downto 0);
    initFilter_return_data : in   std_logic_vector(1 downto 0);
    initFilter_return_tag :  in   std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_call_reqs : out  std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_call_acks : in   std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_call_data : out  std_logic_vector(6 downto 0);
    cal_col_to_be_replaced_call_tag  :  out  std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_return_reqs : out  std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_return_acks : in   std_logic_vector(0 downto 0);
    cal_col_to_be_replaced_return_data : in   std_logic_vector(1 downto 0);
    cal_col_to_be_replaced_return_tag :  in   std_logic_vector(0 downto 0);
    mainAcc_call_reqs : out  std_logic_vector(0 downto 0);
    mainAcc_call_acks : in   std_logic_vector(0 downto 0);
    mainAcc_call_data : out  std_logic_vector(12 downto 0);
    mainAcc_call_tag  :  out  std_logic_vector(0 downto 0);
    mainAcc_return_reqs : out  std_logic_vector(0 downto 0);
    mainAcc_return_acks : in   std_logic_vector(0 downto 0);
    mainAcc_return_data : in   std_logic_vector(15 downto 0);
    mainAcc_return_tag :  in   std_logic_vector(0 downto 0);
    mainAcc2_call_reqs : out  std_logic_vector(0 downto 0);
    mainAcc2_call_acks : in   std_logic_vector(0 downto 0);
    mainAcc2_call_data : out  std_logic_vector(12 downto 0);
    mainAcc2_call_tag  :  out  std_logic_vector(0 downto 0);
    mainAcc2_return_reqs : out  std_logic_vector(0 downto 0);
    mainAcc2_return_acks : in   std_logic_vector(0 downto 0);
    mainAcc2_return_data : in   std_logic_vector(15 downto 0);
    mainAcc2_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accelerator;
architecture accelerator_arch of accelerator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal accelerator_CP_6730_start: Boolean;
  signal accelerator_CP_6730_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component initIfMaps is -- 
    generic (tag_length : integer); 
    port ( -- 
      start : in  std_logic_vector(0 downto 0);
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      finished : out  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component initFilter is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_row_filter : in  std_logic_vector(5 downto 0);
      filter_initialized : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component cal_col_to_be_replaced is -- 
    generic (tag_length : integer); 
    port ( -- 
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      new_col_to_be_replaced : out  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component mainAcc is -- 
    generic (tag_length : integer); 
    port ( -- 
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      ofmap_pixel : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component mainAcc2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      ofmap_pixel : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_1284_ack_0 : boolean;
  signal phi_stmt_1284_req_1 : boolean;
  signal n_I_1335_1288_buf_ack_0 : boolean;
  signal phi_stmt_1284_req_0 : boolean;
  signal n_J_1324_1283_buf_req_1 : boolean;
  signal n_J_1324_1283_buf_req_0 : boolean;
  signal n_J_1324_1283_buf_ack_0 : boolean;
  signal n_I_1335_1288_buf_req_1 : boolean;
  signal n_I_1335_1288_buf_ack_1 : boolean;
  signal n_I_1335_1288_buf_req_0 : boolean;
  signal n_J_1324_1283_buf_ack_1 : boolean;
  signal RPIPE_start_accelerator_1246_inst_req_0 : boolean;
  signal RPIPE_start_accelerator_1246_inst_ack_0 : boolean;
  signal RPIPE_start_accelerator_1246_inst_req_1 : boolean;
  signal RPIPE_start_accelerator_1246_inst_ack_1 : boolean;
  signal if_stmt_1248_branch_req_0 : boolean;
  signal if_stmt_1248_branch_ack_1 : boolean;
  signal if_stmt_1248_branch_ack_0 : boolean;
  signal call_stmt_1259_call_req_0 : boolean;
  signal call_stmt_1259_call_ack_0 : boolean;
  signal call_stmt_1259_call_req_1 : boolean;
  signal call_stmt_1259_call_ack_1 : boolean;
  signal if_stmt_1266_branch_req_0 : boolean;
  signal if_stmt_1266_branch_ack_1 : boolean;
  signal if_stmt_1266_branch_ack_0 : boolean;
  signal do_while_stmt_1271_branch_req_0 : boolean;
  signal phi_stmt_1273_req_1 : boolean;
  signal phi_stmt_1273_req_0 : boolean;
  signal phi_stmt_1273_ack_0 : boolean;
  signal n_ele_1313_1278_buf_req_0 : boolean;
  signal n_ele_1313_1278_buf_ack_0 : boolean;
  signal n_ele_1313_1278_buf_req_1 : boolean;
  signal n_ele_1313_1278_buf_ack_1 : boolean;
  signal phi_stmt_1279_req_1 : boolean;
  signal phi_stmt_1279_req_0 : boolean;
  signal phi_stmt_1279_ack_0 : boolean;
  signal phi_stmt_1289_req_1 : boolean;
  signal phi_stmt_1289_req_0 : boolean;
  signal phi_stmt_1289_ack_0 : boolean;
  signal n_col_to_be_replaced_1342_1293_buf_req_0 : boolean;
  signal n_col_to_be_replaced_1342_1293_buf_ack_0 : boolean;
  signal n_col_to_be_replaced_1342_1293_buf_req_1 : boolean;
  signal n_col_to_be_replaced_1342_1293_buf_ack_1 : boolean;
  signal call_stmt_1307_call_req_0 : boolean;
  signal call_stmt_1307_call_ack_0 : boolean;
  signal call_stmt_1307_call_req_1 : boolean;
  signal call_stmt_1307_call_ack_1 : boolean;
  signal call_stmt_1339_call_req_0 : boolean;
  signal call_stmt_1339_call_ack_0 : boolean;
  signal call_stmt_1339_call_req_1 : boolean;
  signal call_stmt_1339_call_ack_1 : boolean;
  signal call_stmt_1347_call_req_0 : boolean;
  signal call_stmt_1347_call_ack_0 : boolean;
  signal call_stmt_1347_call_req_1 : boolean;
  signal call_stmt_1347_call_ack_1 : boolean;
  signal call_stmt_1363_call_req_0 : boolean;
  signal call_stmt_1363_call_ack_0 : boolean;
  signal call_stmt_1363_call_req_1 : boolean;
  signal call_stmt_1363_call_ack_1 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal WPIPE_read_sums_1364_inst_req_0 : boolean;
  signal WPIPE_read_sums_1364_inst_ack_0 : boolean;
  signal WPIPE_read_sums_1364_inst_req_1 : boolean;
  signal WPIPE_read_sums_1364_inst_ack_1 : boolean;
  signal W_I_1457_delayed_4_0_1368_inst_req_0 : boolean;
  signal W_I_1457_delayed_4_0_1368_inst_ack_0 : boolean;
  signal W_I_1457_delayed_4_0_1368_inst_req_1 : boolean;
  signal W_I_1457_delayed_4_0_1368_inst_ack_1 : boolean;
  signal W_J_1458_delayed_4_0_1371_inst_req_0 : boolean;
  signal W_J_1458_delayed_4_0_1371_inst_ack_0 : boolean;
  signal W_J_1458_delayed_4_0_1371_inst_req_1 : boolean;
  signal W_J_1458_delayed_4_0_1371_inst_ack_1 : boolean;
  signal call_stmt_1379_call_req_0 : boolean;
  signal call_stmt_1379_call_ack_0 : boolean;
  signal call_stmt_1379_call_req_1 : boolean;
  signal call_stmt_1379_call_ack_1 : boolean;
  signal W_checkIFour_1462_delayed_4_0_1380_inst_req_0 : boolean;
  signal W_checkIFour_1462_delayed_4_0_1380_inst_ack_0 : boolean;
  signal W_checkIFour_1462_delayed_4_0_1380_inst_req_1 : boolean;
  signal W_checkIFour_1462_delayed_4_0_1380_inst_ack_1 : boolean;
  signal W_I_1_1464_delayed_4_0_1383_inst_req_0 : boolean;
  signal W_I_1_1464_delayed_4_0_1383_inst_ack_0 : boolean;
  signal W_I_1_1464_delayed_4_0_1383_inst_req_1 : boolean;
  signal W_I_1_1464_delayed_4_0_1383_inst_ack_1 : boolean;
  signal W_J_1465_delayed_4_0_1386_inst_req_0 : boolean;
  signal W_J_1465_delayed_4_0_1386_inst_ack_0 : boolean;
  signal W_J_1465_delayed_4_0_1386_inst_req_1 : boolean;
  signal W_J_1465_delayed_4_0_1386_inst_ack_1 : boolean;
  signal call_stmt_1395_call_req_0 : boolean;
  signal call_stmt_1395_call_ack_0 : boolean;
  signal call_stmt_1395_call_req_1 : boolean;
  signal call_stmt_1395_call_ack_1 : boolean;
  signal do_while_stmt_1271_branch_ack_0 : boolean;
  signal do_while_stmt_1271_branch_ack_1 : boolean;
  signal WPIPE_accelerator_done_1401_inst_req_0 : boolean;
  signal WPIPE_accelerator_done_1401_inst_ack_0 : boolean;
  signal WPIPE_accelerator_done_1401_inst_req_1 : boolean;
  signal WPIPE_accelerator_done_1401_inst_ack_1 : boolean;
  signal phi_stmt_1239_req_0 : boolean;
  signal n_iter_1256_1243_buf_req_0 : boolean;
  signal n_iter_1256_1243_buf_ack_0 : boolean;
  signal n_iter_1256_1243_buf_req_1 : boolean;
  signal n_iter_1256_1243_buf_ack_1 : boolean;
  signal phi_stmt_1239_req_1 : boolean;
  signal phi_stmt_1239_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accelerator_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accelerator_CP_6730_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accelerator_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accelerator_CP_6730_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accelerator_CP_6730_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accelerator_CP_6730_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accelerator_CP_6730_start,"accelerator cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accelerator_CP_6730_symbol, "accelerator cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accelerator_CP_6730: Block -- control-path 
    signal accelerator_CP_6730_elements: BooleanArray(167 downto 0);
    -- 
  begin -- 
    accelerator_CP_6730_elements(0) <= accelerator_CP_6730_start;
    accelerator_CP_6730_symbol <= accelerator_CP_6730_elements(4);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	162 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1237/$entry
      -- CP-element group 0: 	 branch_block_stmt_1237/branch_block_stmt_1237__entry__
      -- CP-element group 0: 	 branch_block_stmt_1237/merge_stmt_1238__entry__
      -- CP-element group 0: 	 branch_block_stmt_1237/merge_stmt_1238_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/$entry
      -- CP-element group 0: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/phi_stmt_1239_sources/$entry
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	167 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Update/cr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:RPIPE_start_accelerator_1246_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:RPIPE_start_accelerator_1246_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_6755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_accelerator_1246_inst_ack_0, ack => accelerator_CP_6730_elements(1)); -- 
    cr_6759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(1), ack => RPIPE_start_accelerator_1246_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_1237/assign_stmt_1247__exit__
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248__entry__
      -- CP-element group 2: 	 branch_block_stmt_1237/assign_stmt_1247/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/EQ_u16_u1_1251_inputs/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/EQ_u16_u1_1251_inputs/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/EQ_u16_u1_1251/SplitProtocol/Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_1237/EQ_u16_u1_1251_place
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1237/if_stmt_1248_else_link/$entry
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:RPIPE_start_accelerator_1246_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1248_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_6760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_start_accelerator_1246_inst_ack_1, ack => accelerator_CP_6730_elements(2)); -- 
    branch_req_6787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(2), ack => if_stmt_1248_branch_req_0); -- 
    -- CP-element group 3:  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	5 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (10) 
      -- CP-element group 3: 	 branch_block_stmt_1237/if_stmt_1248_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_1237/if_stmt_1248_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263__entry__
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/$entry
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1248_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1259_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1259_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_6792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1248_branch_ack_1, ack => accelerator_CP_6730_elements(3)); -- 
    crr_6812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(3), ack => call_stmt_1259_call_req_0); -- 
    ccr_6817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(3), ack => call_stmt_1259_call_req_1); -- 
    -- CP-element group 4:  merge  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 branch_block_stmt_1237/$exit
      -- CP-element group 4: 	 branch_block_stmt_1237/branch_block_stmt_1237__exit__
      -- CP-element group 4: 	 branch_block_stmt_1237/if_stmt_1248__exit__
      -- CP-element group 4: 	 branch_block_stmt_1237/if_stmt_1248_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_1237/if_stmt_1248_else_link/else_choice_transition
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1248_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_6796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1248_branch_ack_0, ack => accelerator_CP_6730_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	3 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1259_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1259_call_ack_0, ack => accelerator_CP_6730_elements(5)); -- 
    -- CP-element group 6:  branch  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	161 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263__exit__
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264__entry__
      -- CP-element group 6: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/$exit
      -- CP-element group 6: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1237/assign_stmt_1256_to_assign_stmt_1263/call_stmt_1259_Update/cca
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/$entry
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1264__entry__
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265__entry__
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265_dead_link/$entry
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265__entry___PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265__entry___PhiReq/$exit
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1259_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_6818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1259_call_ack_1, ack => accelerator_CP_6730_elements(6)); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	161 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_if_link/$exit
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_if_link/if_choice_transition
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270__entry__
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/$entry
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/branch_block_stmt_1270__entry__
      -- CP-element group 7: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271__entry__
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1266_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_6859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1266_branch_ack_1, ack => accelerator_CP_6730_elements(7)); -- 
    -- CP-element group 8:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	161 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	164 
    -- CP-element group 8:  members (15) 
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264__exit__
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264/$exit
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1264__exit__
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266__exit__
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_else_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_else_link/else_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Sample/req
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1266_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_iter_1256_1243_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_iter_1256_1243_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1266_branch_ack_0, ack => accelerator_CP_6730_elements(8)); -- 
    req_7333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(8), ack => n_iter_1256_1243_buf_req_0); -- 
    req_7338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(8), ack => n_iter_1256_1243_buf_req_1); -- 
    -- CP-element group 9:  transition  place  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	158 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	159 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270__exit__
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404__entry__
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/$exit
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/branch_block_stmt_1270__exit__
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271__exit__
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/$entry
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_accelerator_done_1401_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(9), ack => WPIPE_accelerator_done_1401_inst_req_0); -- 
    accelerator_CP_6730_elements(9) <= accelerator_CP_6730_elements(158);
    -- CP-element group 10:  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/$entry
      -- CP-element group 10: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271__entry__
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(10) <= accelerator_CP_6730_elements(7);
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	158 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271__exit__
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(11) is bound as output of CP function.
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_back
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(12) is bound as output of CP function.
    -- CP-element group 13:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	156 
    -- CP-element group 13: 	157 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/condition_done
      -- CP-element group 13: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_exit/$entry
      -- CP-element group 13: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_taken/$entry
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(13) <= accelerator_CP_6730_elements(18);
    -- CP-element group 14:  branch  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	155 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_body_done
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(14) <= accelerator_CP_6730_elements(155);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	46 
    -- CP-element group 15: 	65 
    -- CP-element group 15: 	84 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(15) <= accelerator_CP_6730_elements(12);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16: 	48 
    -- CP-element group 16: 	67 
    -- CP-element group 16: 	86 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(16) <= accelerator_CP_6730_elements(10);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	41 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	60 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	79 
    -- CP-element group 17: 	148 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/$entry
      -- CP-element group 17: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/loop_body_start
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(17) is bound as output of CP function.
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: 	26 
    -- CP-element group 18: 	148 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/condition_evaluated
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:do_while_stmt_1271_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_6890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(18), ack => do_while_stmt_1271_branch_req_0); -- 
    accelerator_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 20,1 => 20,2 => 20);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(22) & accelerator_CP_6730_elements(26) & accelerator_CP_6730_elements(148);
      gj_accelerator_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	40 
    -- CP-element group 19: 	59 
    -- CP-element group 19: 	78 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19: 	80 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/aggregated_phi_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_sample_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 20,1 => 20,2 => 20,3 => 20,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(23) & accelerator_CP_6730_elements(40) & accelerator_CP_6730_elements(59) & accelerator_CP_6730_elements(78) & accelerator_CP_6730_elements(22);
      gj_accelerator_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	62 
    -- CP-element group 20: 	81 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	155 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: 	40 
    -- CP-element group 20: 	59 
    -- CP-element group 20: 	78 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/aggregated_phi_sample_ack
      -- CP-element group 20: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_sample_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 20,1 => 20,2 => 20,3 => 20);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(25) & accelerator_CP_6730_elements(43) & accelerator_CP_6730_elements(62) & accelerator_CP_6730_elements(81);
      gj_accelerator_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21: 	60 
    -- CP-element group 21: 	79 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	44 
    -- CP-element group 21: 	63 
    -- CP-element group 21: 	82 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/aggregated_phi_update_req
      -- CP-element group 21: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_update_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 20,1 => 20,2 => 20,3 => 20);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(24) & accelerator_CP_6730_elements(41) & accelerator_CP_6730_elements(60) & accelerator_CP_6730_elements(79);
      gj_accelerator_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: 	45 
    -- CP-element group 22: 	64 
    -- CP-element group 22: 	83 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 20,1 => 20,2 => 20,3 => 20);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(26) & accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(83);
      gj_accelerator_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	20 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(20);
      gj_accelerator_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	115 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	21 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 20,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(26) & accelerator_CP_6730_elements(115);
      gj_accelerator_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	20 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_sample_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	18 
    -- CP-element group 26: 	22 
    -- CP-element group 26: 	113 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_loopback_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(27) <= accelerator_CP_6730_elements(15);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_loopback_sample_req
      -- CP-element group 28: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_loopback_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1273_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1273_loopback_sample_req_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1273_loopback_sample_req_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(28), ack => phi_stmt_1273_req_1); -- 
    -- Element group accelerator_CP_6730_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_entry_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(29) <= accelerator_CP_6730_elements(16);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_entry_sample_req
      -- CP-element group 30: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_entry_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1273_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1273_entry_sample_req_6908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1273_entry_sample_req_6908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(30), ack => phi_stmt_1273_req_0); -- 
    -- Element group accelerator_CP_6730_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_phi_mux_ack
      -- CP-element group 31: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1273_phi_mux_ack_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1273_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1273_phi_mux_ack_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1273_ack_0, ack => accelerator_CP_6730_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_sample_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(34) <= accelerator_CP_6730_elements(35);
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1277_update_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(33), ack => accelerator_CP_6730_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_sample_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_ele_1313_1278_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_6932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(36), ack => n_ele_1313_1278_buf_req_0); -- 
    -- Element group accelerator_CP_6730_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_update_start__ps
      -- CP-element group 37: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_ele_1313_1278_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_6937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(37), ack => n_ele_1313_1278_buf_req_1); -- 
    -- Element group accelerator_CP_6730_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_ele_1313_1278_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_ele_1313_1278_buf_ack_0, ack => accelerator_CP_6730_elements(38)); -- 
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_ele_1278_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_ele_1313_1278_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_6938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_ele_1313_1278_buf_ack_1, ack => accelerator_CP_6730_elements(39)); -- 
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	20 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	19 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(20);
      gj_accelerator_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	17 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	45 
    -- CP-element group 41: 	99 
    -- CP-element group 41: 	103 
    -- CP-element group 41: 	107 
    -- CP-element group 41: 	111 
    -- CP-element group 41: 	126 
    -- CP-element group 41: 	142 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	21 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 20,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(99) & accelerator_CP_6730_elements(103) & accelerator_CP_6730_elements(107) & accelerator_CP_6730_elements(111) & accelerator_CP_6730_elements(126) & accelerator_CP_6730_elements(142);
      gj_accelerator_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_sample_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(42) <= accelerator_CP_6730_elements(19);
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_sample_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	21 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_update_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(44) <= accelerator_CP_6730_elements(21);
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: 	97 
    -- CP-element group 45: 	101 
    -- CP-element group 45: 	105 
    -- CP-element group 45: 	109 
    -- CP-element group 45: 	124 
    -- CP-element group 45: 	140 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	41 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	15 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_loopback_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(46) <= accelerator_CP_6730_elements(15);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_loopback_sample_req
      -- CP-element group 47: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_loopback_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1279_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1279_loopback_sample_req_6949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1279_loopback_sample_req_6949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(47), ack => phi_stmt_1279_req_1); -- 
    -- Element group accelerator_CP_6730_elements(47) is bound as output of CP function.
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	16 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_entry_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(48) <= accelerator_CP_6730_elements(16);
    -- CP-element group 49:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_entry_sample_req
      -- CP-element group 49: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_entry_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1279_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1279_entry_sample_req_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1279_entry_sample_req_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(49), ack => phi_stmt_1279_req_0); -- 
    -- Element group accelerator_CP_6730_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_phi_mux_ack
      -- CP-element group 50: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1279_phi_mux_ack_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1279_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1279_phi_mux_ack_6955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1279_ack_0, ack => accelerator_CP_6730_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_sample_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_update_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(52) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(53) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(53) <= accelerator_CP_6730_elements(54);
    -- CP-element group 54:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	53 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1282_update_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(54) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(52), ack => accelerator_CP_6730_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_J_1324_1283_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_6976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(55), ack => n_J_1324_1283_buf_req_0); -- 
    -- Element group accelerator_CP_6730_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Update/req
      -- CP-element group 56: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Update/$entry
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_J_1324_1283_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_6981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(56), ack => n_J_1324_1283_buf_req_1); -- 
    -- Element group accelerator_CP_6730_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_J_1324_1283_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_J_1324_1283_buf_ack_0, ack => accelerator_CP_6730_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_J_1283_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_J_1324_1283_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_J_1324_1283_buf_ack_1, ack => accelerator_CP_6730_elements(58)); -- 
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	17 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	20 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	19 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(20);
      gj_accelerator_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	17 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	99 
    -- CP-element group 60: 	107 
    -- CP-element group 60: 	111 
    -- CP-element group 60: 	122 
    -- CP-element group 60: 	134 
    -- CP-element group 60: 	138 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	21 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(60) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 20,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(99) & accelerator_CP_6730_elements(107) & accelerator_CP_6730_elements(111) & accelerator_CP_6730_elements(122) & accelerator_CP_6730_elements(134) & accelerator_CP_6730_elements(138);
      gj_accelerator_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_sample_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(61) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(61) <= accelerator_CP_6730_elements(19);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	20 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_sample_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	21 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_update_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(63) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(63) <= accelerator_CP_6730_elements(21);
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	22 
    -- CP-element group 64: 	97 
    -- CP-element group 64: 	105 
    -- CP-element group 64: 	109 
    -- CP-element group 64: 	120 
    -- CP-element group 64: 	132 
    -- CP-element group 64: 	136 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	15 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_loopback_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(65) <= accelerator_CP_6730_elements(15);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_loopback_sample_req_ps
      -- CP-element group 66: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_loopback_sample_req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1284_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1284_loopback_sample_req_6993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1284_loopback_sample_req_6993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(66), ack => phi_stmt_1284_req_1); -- 
    -- Element group accelerator_CP_6730_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	16 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_entry_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(67) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(67) <= accelerator_CP_6730_elements(16);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_entry_sample_req_ps
      -- CP-element group 68: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_entry_sample_req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1284_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1284_entry_sample_req_6996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1284_entry_sample_req_6996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(68), ack => phi_stmt_1284_req_0); -- 
    -- Element group accelerator_CP_6730_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_phi_mux_ack
      -- CP-element group 69: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1284_phi_mux_ack_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1284_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1284_phi_mux_ack_6999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1284_ack_0, ack => accelerator_CP_6730_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_update_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(72) <= accelerator_CP_6730_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1287_update_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(71), ack => accelerator_CP_6730_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_sample_start__ps
      -- CP-element group 74: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Sample/req
      -- CP-element group 74: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_I_1335_1288_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(74), ack => n_I_1335_1288_buf_req_0); -- 
    -- Element group accelerator_CP_6730_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_update_start__ps
      -- CP-element group 75: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_I_1335_1288_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(75), ack => n_I_1335_1288_buf_req_1); -- 
    -- Element group accelerator_CP_6730_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_I_1335_1288_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_I_1335_1288_buf_ack_0, ack => accelerator_CP_6730_elements(76)); -- 
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_I_1288_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_I_1335_1288_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_I_1335_1288_buf_ack_1, ack => accelerator_CP_6730_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	17 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	20 
    -- CP-element group 78: 	104 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	19 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_sample_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 20,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(20) & accelerator_CP_6730_elements(104);
      gj_accelerator_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	17 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	99 
    -- CP-element group 79: 	103 
    -- CP-element group 79: 	107 
    -- CP-element group 79: 	111 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	21 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(79) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 20,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(17) & accelerator_CP_6730_elements(83) & accelerator_CP_6730_elements(99) & accelerator_CP_6730_elements(103) & accelerator_CP_6730_elements(107) & accelerator_CP_6730_elements(111);
      gj_accelerator_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	19 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_sample_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(80) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(80) <= accelerator_CP_6730_elements(19);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	20 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_sample_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	21 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_update_start__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(82) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(82) <= accelerator_CP_6730_elements(21);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	22 
    -- CP-element group 83: 	97 
    -- CP-element group 83: 	101 
    -- CP-element group 83: 	105 
    -- CP-element group 83: 	109 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(83) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	15 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_loopback_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(84) <= accelerator_CP_6730_elements(15);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_loopback_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_loopback_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1289_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1289_loopback_sample_req_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_loopback_sample_req_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(85), ack => phi_stmt_1289_req_1); -- 
    -- Element group accelerator_CP_6730_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	16 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_entry_trigger
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(86) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(86) <= accelerator_CP_6730_elements(16);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_entry_sample_req
      -- CP-element group 87: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_entry_sample_req_ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1289_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1289_entry_sample_req_7040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_entry_sample_req_7040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(87), ack => phi_stmt_1289_req_0); -- 
    -- Element group accelerator_CP_6730_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_phi_mux_ack_ps
      -- CP-element group 88: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/phi_stmt_1289_phi_mux_ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1289_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1289_phi_mux_ack_7043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1289_ack_0, ack => accelerator_CP_6730_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_sample_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(89) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_update_start_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(90) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_update_completed__ps
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(91) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(91) <= accelerator_CP_6730_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1292_update_completed_
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(92) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(90), ack => accelerator_CP_6730_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_col_to_be_replaced_1342_1293_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(93), ack => n_col_to_be_replaced_1342_1293_buf_req_0); -- 
    -- Element group accelerator_CP_6730_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_col_to_be_replaced_1342_1293_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(94), ack => n_col_to_be_replaced_1342_1293_buf_req_1); -- 
    -- Element group accelerator_CP_6730_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_col_to_be_replaced_1342_1293_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_to_be_replaced_1342_1293_buf_ack_0, ack => accelerator_CP_6730_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/R_n_col_to_be_replaced_1293_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_col_to_be_replaced_1342_1293_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_to_be_replaced_1342_1293_buf_ack_1, ack => accelerator_CP_6730_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	45 
    -- CP-element group 97: 	64 
    -- CP-element group 97: 	83 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	147 
    -- CP-element group 97: 	150 
    -- CP-element group 97: 	154 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1307_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(97), ack => call_stmt_1307_call_req_0); -- 
    accelerator_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 20,1 => 20,2 => 20,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(83) & accelerator_CP_6730_elements(99) & accelerator_CP_6730_elements(147) & accelerator_CP_6730_elements(150) & accelerator_CP_6730_elements(154);
      gj_accelerator_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	100 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1307_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(98), ack => call_stmt_1307_call_req_1); -- 
    accelerator_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accelerator_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accelerator_CP_6730_elements(100);
      gj_accelerator_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	41 
    -- CP-element group 99: 	60 
    -- CP-element group 99: 	79 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1307_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1307_call_ack_0, ack => accelerator_CP_6730_elements(99)); -- 
    -- CP-element group 100:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	149 
    -- CP-element group 100: 	150 
    -- CP-element group 100: 	151 
    -- CP-element group 100: 	153 
    -- CP-element group 100: 	154 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	98 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_Update/cca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1307_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1307_call_ack_1, ack => accelerator_CP_6730_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	45 
    -- CP-element group 101: 	83 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1339_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(101), ack => call_stmt_1339_call_req_0); -- 
    accelerator_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 20,1 => 20,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(83) & accelerator_CP_6730_elements(103);
      gj_accelerator_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1339_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(102), ack => call_stmt_1339_call_req_1); -- 
    accelerator_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(20) & accelerator_CP_6730_elements(104);
      gj_accelerator_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	41 
    -- CP-element group 103: 	79 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1339_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1339_call_ack_0, ack => accelerator_CP_6730_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	155 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	78 
    -- CP-element group 104: 	102 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1339_Update/cca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1339_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1339_call_ack_1, ack => accelerator_CP_6730_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	45 
    -- CP-element group 105: 	64 
    -- CP-element group 105: 	83 
    -- CP-element group 105: 	153 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1347_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(105), ack => call_stmt_1347_call_req_0); -- 
    accelerator_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 20,1 => 20,2 => 20,3 => 20,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(83) & accelerator_CP_6730_elements(153) & accelerator_CP_6730_elements(107);
      gj_accelerator_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: 	130 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1347_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(106), ack => call_stmt_1347_call_req_1); -- 
    accelerator_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(108) & accelerator_CP_6730_elements(130);
      gj_accelerator_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	41 
    -- CP-element group 107: 	60 
    -- CP-element group 107: 	79 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1347_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1347_call_ack_0, ack => accelerator_CP_6730_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	128 
    -- CP-element group 108: 	154 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1347_Update/cca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1347_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1347_call_ack_1, ack => accelerator_CP_6730_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	45 
    -- CP-element group 109: 	64 
    -- CP-element group 109: 	83 
    -- CP-element group 109: 	149 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1363_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(109), ack => call_stmt_1363_call_req_0); -- 
    accelerator_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 20,1 => 20,2 => 20,3 => 20,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(83) & accelerator_CP_6730_elements(149) & accelerator_CP_6730_elements(111);
      gj_accelerator_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: 	146 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1363_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(110), ack => call_stmt_1363_call_req_1); -- 
    accelerator_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(112) & accelerator_CP_6730_elements(146);
      gj_accelerator_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	41 
    -- CP-element group 111: 	60 
    -- CP-element group 111: 	79 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1363_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_0, ack => accelerator_CP_6730_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	144 
    -- CP-element group 112: 	150 
    -- CP-element group 112: 	154 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1363_Update/cca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1363_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_1, ack => accelerator_CP_6730_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	26 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Sample/rr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:type_cast_1366_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(113), ack => type_cast_1366_inst_req_0); -- 
    accelerator_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(26) & accelerator_CP_6730_elements(115);
      gj_accelerator_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: 	118 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_update_start_
      -- CP-element group 114: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Update/cr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:type_cast_1366_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(114), ack => type_cast_1366_inst_req_1); -- 
    accelerator_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(116) & accelerator_CP_6730_elements(118);
      gj_accelerator_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	24 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Sample/ra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:type_cast_1366_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_7136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => accelerator_CP_6730_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/type_cast_1366_Update/ca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:type_cast_1366_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => accelerator_CP_6730_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_read_sums_1364_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(117), ack => WPIPE_read_sums_1364_inst_req_0); -- 
    accelerator_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(116) & accelerator_CP_6730_elements(119);
      gj_accelerator_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	114 
    -- CP-element group 118:  members (6) 
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_update_start_
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Sample/ack
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_read_sums_1364_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_read_sums_1364_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_read_sums_1364_inst_ack_0, ack => accelerator_CP_6730_elements(118)); -- 
    req_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(118), ack => WPIPE_read_sums_1364_inst_req_1); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/WPIPE_read_sums_1364_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_read_sums_1364_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_read_sums_1364_inst_ack_1, ack => accelerator_CP_6730_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	64 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1457_delayed_4_0_1368_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(120), ack => W_I_1457_delayed_4_0_1368_inst_req_0); -- 
    accelerator_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(122);
      gj_accelerator_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	130 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1457_delayed_4_0_1368_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(121), ack => W_I_1457_delayed_4_0_1368_inst_req_1); -- 
    accelerator_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(123) & accelerator_CP_6730_elements(130);
      gj_accelerator_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	60 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1457_delayed_4_0_1368_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_1457_delayed_4_0_1368_inst_ack_0, ack => accelerator_CP_6730_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	128 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1370_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1457_delayed_4_0_1368_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_1457_delayed_4_0_1368_inst_ack_1, ack => accelerator_CP_6730_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	45 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1458_delayed_4_0_1371_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(124), ack => W_J_1458_delayed_4_0_1371_inst_req_0); -- 
    accelerator_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(126);
      gj_accelerator_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	130 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_update_start_
      -- CP-element group 125: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1458_delayed_4_0_1371_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(125), ack => W_J_1458_delayed_4_0_1371_inst_req_1); -- 
    accelerator_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(127) & accelerator_CP_6730_elements(130);
      gj_accelerator_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	41 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1458_delayed_4_0_1371_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_1458_delayed_4_0_1371_inst_ack_0, ack => accelerator_CP_6730_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1373_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1458_delayed_4_0_1371_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_1458_delayed_4_0_1371_inst_ack_1, ack => accelerator_CP_6730_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	108 
    -- CP-element group 128: 	123 
    -- CP-element group 128: 	127 
    -- CP-element group 128: 	151 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1379_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(128), ack => call_stmt_1379_call_req_0); -- 
    accelerator_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 20,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(108) & accelerator_CP_6730_elements(123) & accelerator_CP_6730_elements(127) & accelerator_CP_6730_elements(151) & accelerator_CP_6730_elements(130);
      gj_accelerator_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1379_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(129), ack => call_stmt_1379_call_req_1); -- 
    accelerator_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accelerator_CP_6730_elements(131);
      gj_accelerator_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	106 
    -- CP-element group 130: 	121 
    -- CP-element group 130: 	125 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1379_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1379_call_ack_0, ack => accelerator_CP_6730_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	152 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_Update/cca
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1379_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1379_call_ack_1, ack => accelerator_CP_6730_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	64 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_checkIFour_1462_delayed_4_0_1380_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(132), ack => W_checkIFour_1462_delayed_4_0_1380_inst_req_0); -- 
    accelerator_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(134);
      gj_accelerator_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	146 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_checkIFour_1462_delayed_4_0_1380_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(133), ack => W_checkIFour_1462_delayed_4_0_1380_inst_req_1); -- 
    accelerator_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(135) & accelerator_CP_6730_elements(146);
      gj_accelerator_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	60 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_checkIFour_1462_delayed_4_0_1380_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_checkIFour_1462_delayed_4_0_1380_inst_ack_0, ack => accelerator_CP_6730_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	144 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1382_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_checkIFour_1462_delayed_4_0_1380_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_checkIFour_1462_delayed_4_0_1380_inst_ack_1, ack => accelerator_CP_6730_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	64 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1_1464_delayed_4_0_1383_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(136), ack => W_I_1_1464_delayed_4_0_1383_inst_req_0); -- 
    accelerator_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(64) & accelerator_CP_6730_elements(138);
      gj_accelerator_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	146 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1_1464_delayed_4_0_1383_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(137), ack => W_I_1_1464_delayed_4_0_1383_inst_req_1); -- 
    accelerator_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(139) & accelerator_CP_6730_elements(146);
      gj_accelerator_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	60 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1_1464_delayed_4_0_1383_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_1_1464_delayed_4_0_1383_inst_ack_0, ack => accelerator_CP_6730_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	144 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1385_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_I_1_1464_delayed_4_0_1383_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_1_1464_delayed_4_0_1383_inst_ack_1, ack => accelerator_CP_6730_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	45 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Sample/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1465_delayed_4_0_1386_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(140), ack => W_J_1465_delayed_4_0_1386_inst_req_0); -- 
    accelerator_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(45) & accelerator_CP_6730_elements(142);
      gj_accelerator_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	146 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_update_start_
      -- CP-element group 141: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1465_delayed_4_0_1386_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_7238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(141), ack => W_J_1465_delayed_4_0_1386_inst_req_1); -- 
    accelerator_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(143) & accelerator_CP_6730_elements(146);
      gj_accelerator_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	41 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1465_delayed_4_0_1386_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_1465_delayed_4_0_1386_inst_ack_0, ack => accelerator_CP_6730_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/assign_stmt_1388_Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:W_J_1465_delayed_4_0_1386_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_1465_delayed_4_0_1386_inst_ack_1, ack => accelerator_CP_6730_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	112 
    -- CP-element group 144: 	135 
    -- CP-element group 144: 	139 
    -- CP-element group 144: 	143 
    -- CP-element group 144: 	152 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Sample/crr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1395_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(144), ack => call_stmt_1395_call_req_0); -- 
    accelerator_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 20,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(112) & accelerator_CP_6730_elements(135) & accelerator_CP_6730_elements(139) & accelerator_CP_6730_elements(143) & accelerator_CP_6730_elements(152) & accelerator_CP_6730_elements(146);
      gj_accelerator_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_update_start_
      -- CP-element group 145: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Update/ccr
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1395_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(145), ack => call_stmt_1395_call_req_1); -- 
    accelerator_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accelerator_CP_6730_elements(147);
      gj_accelerator_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	110 
    -- CP-element group 146: 	133 
    -- CP-element group 146: 	137 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Sample/cra
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1395_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1395_call_ack_0, ack => accelerator_CP_6730_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	155 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	97 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1395_Update/cca
      -- CP-element group 147: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/ring_reenable_memory_space_3
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:call_stmt_1395_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1395_call_ack_1, ack => accelerator_CP_6730_elements(147)); -- 
    -- CP-element group 148:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	17 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	18 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(148) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(148) is a control-delay.
    cp_element_148_delay: control_delay_element  generic map(name => " 148_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(17), ack => accelerator_CP_6730_elements(148), clk => clk, reset =>reset);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	100 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	109 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_call_stmt_1363_delay
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(149) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(100), ack => accelerator_CP_6730_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	100 
    -- CP-element group 150: 	112 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	97 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/ring_reenable_memory_space_2
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(150) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 20);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(100) & accelerator_CP_6730_elements(112);
      gj_accelerator_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	100 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	128 
    -- CP-element group 151:  members (1) 
      -- CP-element group 151: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_call_stmt_1379_delay
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(151) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(151) is a control-delay.
    cp_element_151_delay: control_delay_element  generic map(name => " 151_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(100), ack => accelerator_CP_6730_elements(151), clk => clk, reset =>reset);
    -- CP-element group 152:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	131 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	144 
    -- CP-element group 152:  members (1) 
      -- CP-element group 152: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1379_call_stmt_1395_delay
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(152) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(152) is a control-delay.
    cp_element_152_delay: control_delay_element  generic map(name => " 152_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(131), ack => accelerator_CP_6730_elements(152), clk => clk, reset =>reset);
    -- CP-element group 153:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	100 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	105 
    -- CP-element group 153:  members (1) 
      -- CP-element group 153: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/call_stmt_1307_call_stmt_1347_delay
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(153) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accelerator_CP_6730_elements(153) is a control-delay.
    cp_element_153_delay: control_delay_element  generic map(name => " 153_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(100), ack => accelerator_CP_6730_elements(153), clk => clk, reset =>reset);
    -- CP-element group 154:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	100 
    -- CP-element group 154: 	108 
    -- CP-element group 154: 	112 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	97 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/ring_reenable_memory_space_1
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(154) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 20,1 => 20,2 => 20);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(100) & accelerator_CP_6730_elements(108) & accelerator_CP_6730_elements(112);
      gj_accelerator_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	20 
    -- CP-element group 155: 	104 
    -- CP-element group 155: 	119 
    -- CP-element group 155: 	147 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	14 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/do_while_stmt_1271_loop_body/$exit
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(155) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 20,1 => 20,2 => 20,3 => 20,4 => 20,5 => 20);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(20) & accelerator_CP_6730_elements(104) & accelerator_CP_6730_elements(119) & accelerator_CP_6730_elements(147) & accelerator_CP_6730_elements(150) & accelerator_CP_6730_elements(154);
      gj_accelerator_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	13 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_exit/$exit
      -- CP-element group 156: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_exit/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:do_while_stmt_1271_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1271_branch_ack_0, ack => accelerator_CP_6730_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	13 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (2) 
      -- CP-element group 157: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_taken/$exit
      -- CP-element group 157: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/loop_taken/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:do_while_stmt_1271_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1271_branch_ack_1, ack => accelerator_CP_6730_elements(157)); -- 
    -- CP-element group 158:  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	11 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	9 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1237/branch_block_stmt_1264/branch_block_stmt_1270/do_while_stmt_1271/$exit
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(158) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(158) <= accelerator_CP_6730_elements(11);
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	9 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Sample/ack
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Update/req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_accelerator_done_1401_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_accelerator_done_1401_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accelerator_done_1401_inst_ack_0, ack => accelerator_CP_6730_elements(159)); -- 
    req_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(159), ack => WPIPE_accelerator_done_1401_inst_req_1); -- 
    -- CP-element group 160:  transition  place  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (8) 
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404__exit__
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/check_for_filter
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/$exit
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/assign_stmt_1404/WPIPE_accelerator_done_1401_Update/ack
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/check_for_filter_PhiReq/$entry
      -- CP-element group 160: 	 branch_block_stmt_1237/branch_block_stmt_1264/check_for_filter_PhiReq/$exit
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:WPIPE_accelerator_done_1401_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_accelerator_done_1401_inst_ack_1, ack => accelerator_CP_6730_elements(160)); -- 
    -- CP-element group 161:  merge  branch  transition  place  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	6 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	7 
    -- CP-element group 161: 	8 
    -- CP-element group 161:  members (27) 
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265__exit__
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266__entry__
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_dead_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/EQ_u2_u1_1269_inputs/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/EQ_u2_u1_1269_inputs/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Sample/ra
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Update/cr
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/EQ_u2_u1_1269/SplitProtocol/Update/ca
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_eval_test/branch_req
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/EQ_u2_u1_1269_place
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_if_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/if_stmt_1266_else_link/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265_PhiReqMerge
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265_PhiAck/$entry
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265_PhiAck/$exit
      -- CP-element group 161: 	 branch_block_stmt_1237/branch_block_stmt_1264/merge_stmt_1265_PhiAck/dummy
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:if_stmt_1266_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(161), ack => if_stmt_1266_branch_req_0); -- 
    accelerator_CP_6730_elements(161) <= OrReduce(accelerator_CP_6730_elements(6) & accelerator_CP_6730_elements(160));
    -- CP-element group 162:  transition  output  delay-element  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	0 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	166 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/$exit
      -- CP-element group 162: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/$exit
      -- CP-element group 162: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/phi_stmt_1239_sources/$exit
      -- CP-element group 162: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/phi_stmt_1239_sources/type_cast_1242_konst_delay_trans
      -- CP-element group 162: 	 branch_block_stmt_1237/merge_stmt_1238__entry___PhiReq/phi_stmt_1239/phi_stmt_1239_req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1239_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1239_req_7317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1239_req_7317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(162), ack => phi_stmt_1239_req_0); -- 
    -- Element group accelerator_CP_6730_elements(162) is a control-delay.
    cp_element_162_delay: control_delay_element  generic map(name => " 162_delay", delay_value => 1)  port map(req => accelerator_CP_6730_elements(0), ack => accelerator_CP_6730_elements(162), clk => clk, reset =>reset);
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_iter_1256_1243_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iter_1256_1243_buf_ack_0, ack => accelerator_CP_6730_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	8 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:n_iter_1256_1243_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_iter_1256_1243_buf_ack_1, ack => accelerator_CP_6730_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_1237/check_for_start_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/$exit
      -- CP-element group 165: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/$exit
      -- CP-element group 165: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_sources/Interlock/$exit
      -- CP-element group 165: 	 branch_block_stmt_1237/check_for_start_PhiReq/phi_stmt_1239/phi_stmt_1239_req
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1239_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1239_req_7340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1239_req_7340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(165), ack => phi_stmt_1239_req_1); -- 
    accelerator_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accelerator_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accelerator_CP_6730_elements(163) & accelerator_CP_6730_elements(164);
      gj_accelerator_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accelerator_CP_6730_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  merge  transition  place  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	162 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_1237/merge_stmt_1238_PhiReqMerge
      -- CP-element group 166: 	 branch_block_stmt_1237/merge_stmt_1238_PhiAck/$entry
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(166) fired."); 
        -- 
      end if; --
    end process; 
    accelerator_CP_6730_elements(166) <= OrReduce(accelerator_CP_6730_elements(162) & accelerator_CP_6730_elements(165));
    -- CP-element group 167:  merge  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	1 
    -- CP-element group 167:  members (8) 
      -- CP-element group 167: 	 branch_block_stmt_1237/merge_stmt_1238__exit__
      -- CP-element group 167: 	 branch_block_stmt_1237/assign_stmt_1247__entry__
      -- CP-element group 167: 	 branch_block_stmt_1237/assign_stmt_1247/$entry
      -- CP-element group 167: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_1237/assign_stmt_1247/RPIPE_start_accelerator_1246_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_1237/merge_stmt_1238_PhiAck/$exit
      -- CP-element group 167: 	 branch_block_stmt_1237/merge_stmt_1238_PhiAck/phi_stmt_1239_ack
      -- 
    -- logger for CP element group accelerator_CP_6730_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accelerator_CP_6730_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:accelerator_CP_6730_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:phi_stmt_1239_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accelerator:CP:RPIPE_start_accelerator_1246_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1239_ack_7345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1239_ack_0, ack => accelerator_CP_6730_elements(167)); -- 
    rr_6754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accelerator_CP_6730_elements(167), ack => RPIPE_start_accelerator_1246_inst_req_0); -- 
    accelerator_do_while_stmt_1271_terminator_7270: loop_terminator -- 
      generic map (name => " accelerator_do_while_stmt_1271_terminator_7270", max_iterations_in_flight =>20) 
      port map(loop_body_exit => accelerator_CP_6730_elements(14),loop_continue => accelerator_CP_6730_elements(157),loop_terminate => accelerator_CP_6730_elements(156),loop_back => accelerator_CP_6730_elements(12),loop_exit => accelerator_CP_6730_elements(11),clk => clk, reset => reset); -- 
    phi_stmt_1273_phi_seq_6939_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accelerator_CP_6730_elements(29);
      accelerator_CP_6730_elements(32)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accelerator_CP_6730_elements(32);
      accelerator_CP_6730_elements(33)<= src_update_reqs(0);
      src_update_acks(0)  <= accelerator_CP_6730_elements(34);
      accelerator_CP_6730_elements(30) <= phi_mux_reqs(0);
      triggers(1)  <= accelerator_CP_6730_elements(27);
      accelerator_CP_6730_elements(36)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accelerator_CP_6730_elements(38);
      accelerator_CP_6730_elements(37)<= src_update_reqs(1);
      src_update_acks(1)  <= accelerator_CP_6730_elements(39);
      accelerator_CP_6730_elements(28) <= phi_mux_reqs(1);
      phi_stmt_1273_phi_seq_6939 : phi_sequencer_v2-- 
        generic map (place_capacity => 20, ntriggers => 2, name => "phi_stmt_1273_phi_seq_6939") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accelerator_CP_6730_elements(19), 
          phi_sample_ack => accelerator_CP_6730_elements(25), 
          phi_update_req => accelerator_CP_6730_elements(21), 
          phi_update_ack => accelerator_CP_6730_elements(26), 
          phi_mux_ack => accelerator_CP_6730_elements(31), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1279_phi_seq_6983_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accelerator_CP_6730_elements(48);
      accelerator_CP_6730_elements(51)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accelerator_CP_6730_elements(51);
      accelerator_CP_6730_elements(52)<= src_update_reqs(0);
      src_update_acks(0)  <= accelerator_CP_6730_elements(53);
      accelerator_CP_6730_elements(49) <= phi_mux_reqs(0);
      triggers(1)  <= accelerator_CP_6730_elements(46);
      accelerator_CP_6730_elements(55)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accelerator_CP_6730_elements(57);
      accelerator_CP_6730_elements(56)<= src_update_reqs(1);
      src_update_acks(1)  <= accelerator_CP_6730_elements(58);
      accelerator_CP_6730_elements(47) <= phi_mux_reqs(1);
      phi_stmt_1279_phi_seq_6983 : phi_sequencer_v2-- 
        generic map (place_capacity => 20, ntriggers => 2, name => "phi_stmt_1279_phi_seq_6983") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accelerator_CP_6730_elements(42), 
          phi_sample_ack => accelerator_CP_6730_elements(43), 
          phi_update_req => accelerator_CP_6730_elements(44), 
          phi_update_ack => accelerator_CP_6730_elements(45), 
          phi_mux_ack => accelerator_CP_6730_elements(50), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1284_phi_seq_7027_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accelerator_CP_6730_elements(67);
      accelerator_CP_6730_elements(70)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accelerator_CP_6730_elements(70);
      accelerator_CP_6730_elements(71)<= src_update_reqs(0);
      src_update_acks(0)  <= accelerator_CP_6730_elements(72);
      accelerator_CP_6730_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= accelerator_CP_6730_elements(65);
      accelerator_CP_6730_elements(74)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accelerator_CP_6730_elements(76);
      accelerator_CP_6730_elements(75)<= src_update_reqs(1);
      src_update_acks(1)  <= accelerator_CP_6730_elements(77);
      accelerator_CP_6730_elements(66) <= phi_mux_reqs(1);
      phi_stmt_1284_phi_seq_7027 : phi_sequencer_v2-- 
        generic map (place_capacity => 20, ntriggers => 2, name => "phi_stmt_1284_phi_seq_7027") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accelerator_CP_6730_elements(61), 
          phi_sample_ack => accelerator_CP_6730_elements(62), 
          phi_update_req => accelerator_CP_6730_elements(63), 
          phi_update_ack => accelerator_CP_6730_elements(64), 
          phi_mux_ack => accelerator_CP_6730_elements(69), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1289_phi_seq_7071_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accelerator_CP_6730_elements(86);
      accelerator_CP_6730_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accelerator_CP_6730_elements(89);
      accelerator_CP_6730_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= accelerator_CP_6730_elements(91);
      accelerator_CP_6730_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= accelerator_CP_6730_elements(84);
      accelerator_CP_6730_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accelerator_CP_6730_elements(95);
      accelerator_CP_6730_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= accelerator_CP_6730_elements(96);
      accelerator_CP_6730_elements(85) <= phi_mux_reqs(1);
      phi_stmt_1289_phi_seq_7071 : phi_sequencer_v2-- 
        generic map (place_capacity => 20, ntriggers => 2, name => "phi_stmt_1289_phi_seq_7071") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accelerator_CP_6730_elements(80), 
          phi_sample_ack => accelerator_CP_6730_elements(81), 
          phi_update_req => accelerator_CP_6730_elements(82), 
          phi_update_ack => accelerator_CP_6730_elements(83), 
          phi_mux_ack => accelerator_CP_6730_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6891_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= accelerator_CP_6730_elements(15);
        preds(1)  <= accelerator_CP_6730_elements(16);
        entry_tmerge_6891 : transition_merge -- 
          generic map(name => " entry_tmerge_6891")
          port map (preds => preds, symbol_out => accelerator_CP_6730_elements(17));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_1320_wire : std_logic_vector(4 downto 0);
    signal ADD_u6_u6_1298_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1331_wire : std_logic_vector(5 downto 0);
    signal ADD_u7_u7_1311_wire : std_logic_vector(6 downto 0);
    signal EQ_u16_u1_1251_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1269_wire : std_logic_vector(0 downto 0);
    signal EQ_u5_u1_1328_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1351_wire : std_logic_vector(0 downto 0);
    signal I_1284 : std_logic_vector(5 downto 0);
    signal I_1457_delayed_4_0_1370 : std_logic_vector(5 downto 0);
    signal I_1_1300 : std_logic_vector(5 downto 0);
    signal I_1_1464_delayed_4_0_1385 : std_logic_vector(5 downto 0);
    signal J_1279 : std_logic_vector(4 downto 0);
    signal J_1458_delayed_4_0_1373 : std_logic_vector(4 downto 0);
    signal J_1465_delayed_4_0_1388 : std_logic_vector(4 downto 0);
    signal R_filter_start_addr_1257_wire_constant : std_logic_vector(5 downto 0);
    signal R_write_signal_1374_wire_constant : std_logic_vector(0 downto 0);
    signal R_write_signal_1390_wire_constant : std_logic_vector(0 downto 0);
    signal ULT_u5_u1_1317_wire : std_logic_vector(0 downto 0);
    signal ULT_u7_u1_1399_wire : std_logic_vector(0 downto 0);
    signal checkIFour_1357 : std_logic_vector(0 downto 0);
    signal checkIFour_1462_delayed_4_0_1382 : std_logic_vector(0 downto 0);
    signal check_both_1263 : std_logic_vector(1 downto 0);
    signal cmd_1247 : std_logic_vector(15 downto 0);
    signal col_to_be_replaced_1289 : std_logic_vector(1 downto 0);
    signal ele_1273 : std_logic_vector(6 downto 0);
    signal initialized_filter_1259 : std_logic_vector(1 downto 0);
    signal initialized_ifmaps_1307 : std_logic_vector(1 downto 0);
    signal iter_1239 : std_logic_vector(15 downto 0);
    signal konst_1254_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1268_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1297_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1310_wire_constant : std_logic_vector(6 downto 0);
    signal konst_1316_wire_constant : std_logic_vector(4 downto 0);
    signal konst_1319_wire_constant : std_logic_vector(4 downto 0);
    signal konst_1327_wire_constant : std_logic_vector(4 downto 0);
    signal konst_1330_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1350_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1398_wire_constant : std_logic_vector(6 downto 0);
    signal n_I_1335 : std_logic_vector(5 downto 0);
    signal n_I_1335_1288_buffered : std_logic_vector(5 downto 0);
    signal n_J_1324 : std_logic_vector(4 downto 0);
    signal n_J_1324_1283_buffered : std_logic_vector(4 downto 0);
    signal n_col_to_be_replaced_1342 : std_logic_vector(1 downto 0);
    signal n_col_to_be_replaced_1342_1293_buffered : std_logic_vector(1 downto 0);
    signal n_ele_1313 : std_logic_vector(6 downto 0);
    signal n_ele_1313_1278_buffered : std_logic_vector(6 downto 0);
    signal n_iter_1256 : std_logic_vector(15 downto 0);
    signal n_iter_1256_1243_buffered : std_logic_vector(15 downto 0);
    signal new_col_to_be_replaced_1339 : std_logic_vector(1 downto 0);
    signal ofmap_pixel2_1363 : std_logic_vector(15 downto 0);
    signal ofmap_pixel_1347 : std_logic_vector(15 downto 0);
    signal r_data_sum_cal2_1395 : std_logic_vector(15 downto 0);
    signal r_data_sum_cal_1379 : std_logic_vector(15 downto 0);
    signal type_cast_1242_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1277_wire_constant : std_logic_vector(6 downto 0);
    signal type_cast_1282_wire_constant : std_logic_vector(4 downto 0);
    signal type_cast_1287_wire_constant : std_logic_vector(5 downto 0);
    signal type_cast_1292_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_1302_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(4 downto 0);
    signal type_cast_1332_wire : std_logic_vector(5 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1355_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1366_wire : std_logic_vector(15 downto 0);
    signal type_cast_1403_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_filter_start_addr_1257_wire_constant <= "001000";
    R_write_signal_1374_wire_constant <= "0";
    R_write_signal_1390_wire_constant <= "0";
    konst_1254_wire_constant <= "0000000000000001";
    konst_1268_wire_constant <= "01";
    konst_1297_wire_constant <= "000001";
    konst_1310_wire_constant <= "0000001";
    konst_1316_wire_constant <= "00100";
    konst_1319_wire_constant <= "00001";
    konst_1327_wire_constant <= "00100";
    konst_1330_wire_constant <= "000010";
    konst_1350_wire_constant <= "000100";
    konst_1398_wire_constant <= "0001110";
    type_cast_1242_wire_constant <= "0000000000000001";
    type_cast_1277_wire_constant <= "0000000";
    type_cast_1282_wire_constant <= "00000";
    type_cast_1287_wire_constant <= "000000";
    type_cast_1292_wire_constant <= "11";
    type_cast_1302_wire_constant <= "1";
    type_cast_1322_wire_constant <= "00000";
    type_cast_1353_wire_constant <= "1";
    type_cast_1355_wire_constant <= "0";
    type_cast_1403_wire_constant <= "0000000000000001";
    -- logger for phi phi_stmt_1239
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1239_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1239:input-0 type_cast_1242_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1242_wire_constant));
          --
        end if;
        if phi_stmt_1239_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1239:input-1 n_iter_1256_1243_buffered= " & Convert_SLV_To_Hex_String(n_iter_1256_1243_buffered));
          --
        end if;
        if phi_stmt_1239_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:accelerator:DP:phi_stmt_1239:sample-completed");
          --
        end if;
        if phi_stmt_1239_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:accelerator:DP:phi_stmt_1239:output iter_1239= " & Convert_SLV_To_Hex_String(iter_1239));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1239: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1242_wire_constant & n_iter_1256_1243_buffered;
      req <= phi_stmt_1239_req_0 & phi_stmt_1239_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1239",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1239_ack_0,
          idata => idata,
          odata => iter_1239,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1239
    -- logger for phi phi_stmt_1273
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1273_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1273:input-0 type_cast_1277_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1277_wire_constant));
          --
        end if;
        if phi_stmt_1273_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1273:input-1 n_ele_1313_1278_buffered= " & Convert_SLV_To_Hex_String(n_ele_1313_1278_buffered));
          --
        end if;
        if phi_stmt_1273_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:accelerator:DP:phi_stmt_1273:sample-completed");
          --
        end if;
        if phi_stmt_1273_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:accelerator:DP:phi_stmt_1273:output ele_1273= " & Convert_SLV_To_Hex_String(ele_1273));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1273: Block -- phi operator 
      signal idata: std_logic_vector(13 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1277_wire_constant & n_ele_1313_1278_buffered;
      req <= phi_stmt_1273_req_0 & phi_stmt_1273_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1273",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 7) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1273_ack_0,
          idata => idata,
          odata => ele_1273,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1273
    -- logger for phi phi_stmt_1279
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1279_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1279:input-0 type_cast_1282_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1282_wire_constant));
          --
        end if;
        if phi_stmt_1279_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1279:input-1 n_J_1324_1283_buffered= " & Convert_SLV_To_Hex_String(n_J_1324_1283_buffered));
          --
        end if;
        if phi_stmt_1279_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:accelerator:DP:phi_stmt_1279:sample-completed");
          --
        end if;
        if phi_stmt_1279_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:accelerator:DP:phi_stmt_1279:output J_1279= " & Convert_SLV_To_Hex_String(J_1279));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1279: Block -- phi operator 
      signal idata: std_logic_vector(9 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1282_wire_constant & n_J_1324_1283_buffered;
      req <= phi_stmt_1279_req_0 & phi_stmt_1279_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1279",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 5) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1279_ack_0,
          idata => idata,
          odata => J_1279,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1279
    -- logger for phi phi_stmt_1284
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1284_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1284:input-0 type_cast_1287_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1287_wire_constant));
          --
        end if;
        if phi_stmt_1284_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1284:input-1 n_I_1335_1288_buffered= " & Convert_SLV_To_Hex_String(n_I_1335_1288_buffered));
          --
        end if;
        if phi_stmt_1284_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:accelerator:DP:phi_stmt_1284:sample-completed");
          --
        end if;
        if phi_stmt_1284_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:accelerator:DP:phi_stmt_1284:output I_1284= " & Convert_SLV_To_Hex_String(I_1284));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1284: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1287_wire_constant & n_I_1335_1288_buffered;
      req <= phi_stmt_1284_req_0 & phi_stmt_1284_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1284",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1284_ack_0,
          idata => idata,
          odata => I_1284,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1284
    -- logger for phi phi_stmt_1289
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1289_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1289:input-0 type_cast_1292_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_1292_wire_constant));
          --
        end if;
        if phi_stmt_1289_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:accelerator:DP:phi_stmt_1289:input-1 n_col_to_be_replaced_1342_1293_buffered= " & Convert_SLV_To_Hex_String(n_col_to_be_replaced_1342_1293_buffered));
          --
        end if;
        if phi_stmt_1289_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:accelerator:DP:phi_stmt_1289:sample-completed");
          --
        end if;
        if phi_stmt_1289_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:accelerator:DP:phi_stmt_1289:output col_to_be_replaced_1289= " & Convert_SLV_To_Hex_String(col_to_be_replaced_1289));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1289: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1292_wire_constant & n_col_to_be_replaced_1342_1293_buffered;
      req <= phi_stmt_1289_req_0 & phi_stmt_1289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1289",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1289_ack_0,
          idata => idata,
          odata => col_to_be_replaced_1289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1289
    -- logger for split-operator MUX_1323_inst flow-through 
    process(n_J_1324) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:MUX_1323_inst:flowthrough inputs: " & " ULT_u5_u1_1317_wire = "& Convert_SLV_To_Hex_String(ULT_u5_u1_1317_wire) & " ADD_u5_u5_1320_wire = "& Convert_SLV_To_Hex_String(ADD_u5_u5_1320_wire) & " type_cast_1322_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1322_wire_constant) & " outputs:" & " n_J_1324= "  & Convert_SLV_To_Hex_String(n_J_1324));
      --
    end process; 
    -- flow-through select operator MUX_1323_inst
    n_J_1324 <= ADD_u5_u5_1320_wire when (ULT_u5_u1_1317_wire(0) /=  '0') else type_cast_1322_wire_constant;
    -- logger for split-operator MUX_1334_inst flow-through 
    process(n_I_1335) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:MUX_1334_inst:flowthrough inputs: " & " EQ_u5_u1_1328_wire = "& Convert_SLV_To_Hex_String(EQ_u5_u1_1328_wire) & " type_cast_1332_wire = "& Convert_SLV_To_Hex_String(type_cast_1332_wire) & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " outputs:" & " n_I_1335= "  & Convert_SLV_To_Hex_String(n_I_1335));
      --
    end process; 
    -- flow-through select operator MUX_1334_inst
    n_I_1335 <= type_cast_1332_wire when (EQ_u5_u1_1328_wire(0) /=  '0') else I_1284;
    -- logger for split-operator MUX_1356_inst flow-through 
    process(checkIFour_1357) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:MUX_1356_inst:flowthrough inputs: " & " EQ_u6_u1_1351_wire = "& Convert_SLV_To_Hex_String(EQ_u6_u1_1351_wire) & " type_cast_1353_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1353_wire_constant) & " type_cast_1355_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1355_wire_constant) & " outputs:" & " checkIFour_1357= "  & Convert_SLV_To_Hex_String(checkIFour_1357));
      --
    end process; 
    -- flow-through select operator MUX_1356_inst
    checkIFour_1357 <= type_cast_1353_wire_constant when (EQ_u6_u1_1351_wire(0) /=  '0') else type_cast_1355_wire_constant;
    -- logger for split-operator W_I_1457_delayed_4_0_1368_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_I_1457_delayed_4_0_1368_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_I_1457_delayed_4_0_1368_inst:started:   inputs: " & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284));
          --
        end if; 
        if W_I_1457_delayed_4_0_1368_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_I_1457_delayed_4_0_1368_inst:finished:  outputs: " & " I_1457_delayed_4_0_1370= "  & Convert_SLV_To_Hex_String(I_1457_delayed_4_0_1370));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_I_1457_delayed_4_0_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_I_1457_delayed_4_0_1368_inst_req_0;
      W_I_1457_delayed_4_0_1368_inst_ack_0<= wack(0);
      rreq(0) <= W_I_1457_delayed_4_0_1368_inst_req_1;
      W_I_1457_delayed_4_0_1368_inst_ack_1<= rack(0);
      W_I_1457_delayed_4_0_1368_inst : InterlockBuffer generic map ( -- 
        name => "W_I_1457_delayed_4_0_1368_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_1284,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => I_1457_delayed_4_0_1370,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_I_1_1464_delayed_4_0_1383_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_I_1_1464_delayed_4_0_1383_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_I_1_1464_delayed_4_0_1383_inst:started:   inputs: " & " I_1_1300 = "& Convert_SLV_To_Hex_String(I_1_1300));
          --
        end if; 
        if W_I_1_1464_delayed_4_0_1383_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_I_1_1464_delayed_4_0_1383_inst:finished:  outputs: " & " I_1_1464_delayed_4_0_1385= "  & Convert_SLV_To_Hex_String(I_1_1464_delayed_4_0_1385));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_I_1_1464_delayed_4_0_1383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_I_1_1464_delayed_4_0_1383_inst_req_0;
      W_I_1_1464_delayed_4_0_1383_inst_ack_0<= wack(0);
      rreq(0) <= W_I_1_1464_delayed_4_0_1383_inst_req_1;
      W_I_1_1464_delayed_4_0_1383_inst_ack_1<= rack(0);
      W_I_1_1464_delayed_4_0_1383_inst : InterlockBuffer generic map ( -- 
        name => "W_I_1_1464_delayed_4_0_1383_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_1_1300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => I_1_1464_delayed_4_0_1385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_J_1458_delayed_4_0_1371_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_J_1458_delayed_4_0_1371_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_J_1458_delayed_4_0_1371_inst:started:   inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279));
          --
        end if; 
        if W_J_1458_delayed_4_0_1371_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_J_1458_delayed_4_0_1371_inst:finished:  outputs: " & " J_1458_delayed_4_0_1373= "  & Convert_SLV_To_Hex_String(J_1458_delayed_4_0_1373));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_J_1458_delayed_4_0_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_J_1458_delayed_4_0_1371_inst_req_0;
      W_J_1458_delayed_4_0_1371_inst_ack_0<= wack(0);
      rreq(0) <= W_J_1458_delayed_4_0_1371_inst_req_1;
      W_J_1458_delayed_4_0_1371_inst_ack_1<= rack(0);
      W_J_1458_delayed_4_0_1371_inst : InterlockBuffer generic map ( -- 
        name => "W_J_1458_delayed_4_0_1371_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => J_1279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => J_1458_delayed_4_0_1373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_J_1465_delayed_4_0_1386_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_J_1465_delayed_4_0_1386_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_J_1465_delayed_4_0_1386_inst:started:   inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279));
          --
        end if; 
        if W_J_1465_delayed_4_0_1386_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_J_1465_delayed_4_0_1386_inst:finished:  outputs: " & " J_1465_delayed_4_0_1388= "  & Convert_SLV_To_Hex_String(J_1465_delayed_4_0_1388));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_J_1465_delayed_4_0_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_J_1465_delayed_4_0_1386_inst_req_0;
      W_J_1465_delayed_4_0_1386_inst_ack_0<= wack(0);
      rreq(0) <= W_J_1465_delayed_4_0_1386_inst_req_1;
      W_J_1465_delayed_4_0_1386_inst_ack_1<= rack(0);
      W_J_1465_delayed_4_0_1386_inst : InterlockBuffer generic map ( -- 
        name => "W_J_1465_delayed_4_0_1386_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => J_1279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => J_1465_delayed_4_0_1388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_checkIFour_1462_delayed_4_0_1380_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_checkIFour_1462_delayed_4_0_1380_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_checkIFour_1462_delayed_4_0_1380_inst:started:   inputs: " & " checkIFour_1357 = "& Convert_SLV_To_Hex_String(checkIFour_1357));
          --
        end if; 
        if W_checkIFour_1462_delayed_4_0_1380_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_checkIFour_1462_delayed_4_0_1380_inst:finished:  outputs: " & " checkIFour_1462_delayed_4_0_1382= "  & Convert_SLV_To_Hex_String(checkIFour_1462_delayed_4_0_1382));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_checkIFour_1462_delayed_4_0_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_checkIFour_1462_delayed_4_0_1380_inst_req_0;
      W_checkIFour_1462_delayed_4_0_1380_inst_ack_0<= wack(0);
      rreq(0) <= W_checkIFour_1462_delayed_4_0_1380_inst_req_1;
      W_checkIFour_1462_delayed_4_0_1380_inst_ack_1<= rack(0);
      W_checkIFour_1462_delayed_4_0_1380_inst : InterlockBuffer generic map ( -- 
        name => "W_checkIFour_1462_delayed_4_0_1380_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => checkIFour_1357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => checkIFour_1462_delayed_4_0_1382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_n_col_to_be_replaced_1340_inst flow-through 
    process(n_col_to_be_replaced_1342) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:W_n_col_to_be_replaced_1340_inst:flowthrough inputs: " & " new_col_to_be_replaced_1339 = "& Convert_SLV_To_Hex_String(new_col_to_be_replaced_1339) & " outputs:" & " n_col_to_be_replaced_1342= "  & Convert_SLV_To_Hex_String(n_col_to_be_replaced_1342));
      --
    end process; 
    -- interlock W_n_col_to_be_replaced_1340_inst
    process(new_col_to_be_replaced_1339) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := new_col_to_be_replaced_1339(1 downto 0);
      n_col_to_be_replaced_1342 <= tmp_var; -- 
    end process;
    -- logger for split-operator n_I_1335_1288_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_I_1335_1288_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_I_1335_1288_buf:started:   inputs: " & " n_I_1335 = "& Convert_SLV_To_Hex_String(n_I_1335));
          --
        end if; 
        if n_I_1335_1288_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_I_1335_1288_buf:finished:  outputs: " & " n_I_1335_1288_buffered= "  & Convert_SLV_To_Hex_String(n_I_1335_1288_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_I_1335_1288_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_I_1335_1288_buf_req_0;
      n_I_1335_1288_buf_ack_0<= wack(0);
      rreq(0) <= n_I_1335_1288_buf_req_1;
      n_I_1335_1288_buf_ack_1<= rack(0);
      n_I_1335_1288_buf : InterlockBuffer generic map ( -- 
        name => "n_I_1335_1288_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_I_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_I_1335_1288_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_J_1324_1283_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_J_1324_1283_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_J_1324_1283_buf:started:   inputs: " & " n_J_1324 = "& Convert_SLV_To_Hex_String(n_J_1324));
          --
        end if; 
        if n_J_1324_1283_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_J_1324_1283_buf:finished:  outputs: " & " n_J_1324_1283_buffered= "  & Convert_SLV_To_Hex_String(n_J_1324_1283_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_J_1324_1283_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_J_1324_1283_buf_req_0;
      n_J_1324_1283_buf_ack_0<= wack(0);
      rreq(0) <= n_J_1324_1283_buf_req_1;
      n_J_1324_1283_buf_ack_1<= rack(0);
      n_J_1324_1283_buf : InterlockBuffer generic map ( -- 
        name => "n_J_1324_1283_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_J_1324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_J_1324_1283_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_col_to_be_replaced_1342_1293_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_col_to_be_replaced_1342_1293_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_col_to_be_replaced_1342_1293_buf:started:   inputs: " & " n_col_to_be_replaced_1342 = "& Convert_SLV_To_Hex_String(n_col_to_be_replaced_1342));
          --
        end if; 
        if n_col_to_be_replaced_1342_1293_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_col_to_be_replaced_1342_1293_buf:finished:  outputs: " & " n_col_to_be_replaced_1342_1293_buffered= "  & Convert_SLV_To_Hex_String(n_col_to_be_replaced_1342_1293_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_col_to_be_replaced_1342_1293_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_to_be_replaced_1342_1293_buf_req_0;
      n_col_to_be_replaced_1342_1293_buf_ack_0<= wack(0);
      rreq(0) <= n_col_to_be_replaced_1342_1293_buf_req_1;
      n_col_to_be_replaced_1342_1293_buf_ack_1<= rack(0);
      n_col_to_be_replaced_1342_1293_buf : InterlockBuffer generic map ( -- 
        name => "n_col_to_be_replaced_1342_1293_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_to_be_replaced_1342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_to_be_replaced_1342_1293_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_ele_1313_1278_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_ele_1313_1278_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_ele_1313_1278_buf:started:   inputs: " & " n_ele_1313 = "& Convert_SLV_To_Hex_String(n_ele_1313));
          --
        end if; 
        if n_ele_1313_1278_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_ele_1313_1278_buf:finished:  outputs: " & " n_ele_1313_1278_buffered= "  & Convert_SLV_To_Hex_String(n_ele_1313_1278_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_ele_1313_1278_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_ele_1313_1278_buf_req_0;
      n_ele_1313_1278_buf_ack_0<= wack(0);
      rreq(0) <= n_ele_1313_1278_buf_req_1;
      n_ele_1313_1278_buf_ack_1<= rack(0);
      n_ele_1313_1278_buf : InterlockBuffer generic map ( -- 
        name => "n_ele_1313_1278_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 7,
        out_data_width => 7,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_ele_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_ele_1313_1278_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_iter_1256_1243_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_iter_1256_1243_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_iter_1256_1243_buf:started:   inputs: " & " n_iter_1256 = "& Convert_SLV_To_Hex_String(n_iter_1256));
          --
        end if; 
        if n_iter_1256_1243_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:n_iter_1256_1243_buf:finished:  outputs: " & " n_iter_1256_1243_buffered= "  & Convert_SLV_To_Hex_String(n_iter_1256_1243_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_iter_1256_1243_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_iter_1256_1243_buf_req_0;
      n_iter_1256_1243_buf_ack_0<= wack(0);
      rreq(0) <= n_iter_1256_1243_buf_req_1;
      n_iter_1256_1243_buf_ack_1<= rack(0);
      n_iter_1256_1243_buf : InterlockBuffer generic map ( -- 
        name => "n_iter_1256_1243_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_iter_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_iter_1256_1243_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1262_inst flow-through 
    process(check_both_1263) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1262_inst:flowthrough inputs: " & " initialized_filter_1259 = "& Convert_SLV_To_Hex_String(initialized_filter_1259) & " outputs:" & " check_both_1263= "  & Convert_SLV_To_Hex_String(check_both_1263));
      --
    end process; 
    -- interlock type_cast_1262_inst
    process(initialized_filter_1259) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := initialized_filter_1259(1 downto 0);
      check_both_1263 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1299_inst flow-through 
    process(I_1_1300) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1299_inst:flowthrough inputs: " & " ADD_u6_u6_1298_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_1298_wire) & " outputs:" & " I_1_1300= "  & Convert_SLV_To_Hex_String(I_1_1300));
      --
    end process; 
    -- interlock type_cast_1299_inst
    process(ADD_u6_u6_1298_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1298_wire(5 downto 0);
      I_1_1300 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1312_inst flow-through 
    process(n_ele_1313) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1312_inst:flowthrough inputs: " & " ADD_u7_u7_1311_wire = "& Convert_SLV_To_Hex_String(ADD_u7_u7_1311_wire) & " outputs:" & " n_ele_1313= "  & Convert_SLV_To_Hex_String(n_ele_1313));
      --
    end process; 
    -- interlock type_cast_1312_inst
    process(ADD_u7_u7_1311_wire) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 6 downto 0) := ADD_u7_u7_1311_wire(6 downto 0);
      n_ele_1313 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1332_inst flow-through 
    process(type_cast_1332_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1332_inst:flowthrough inputs: " & " ADD_u6_u6_1331_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_1331_wire) & " outputs:" & " type_cast_1332_wire= "  & Convert_SLV_To_Hex_String(type_cast_1332_wire));
      --
    end process; 
    -- interlock type_cast_1332_inst
    process(ADD_u6_u6_1331_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1331_wire(5 downto 0);
      type_cast_1332_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1366_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1366_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1366_inst:started:   inputs: " & " ele_1273 = "& Convert_SLV_To_Hex_String(ele_1273));
          --
        end if; 
        if type_cast_1366_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:type_cast_1366_inst:finished:  outputs: " & " type_cast_1366_wire= "  & Convert_SLV_To_Hex_String(type_cast_1366_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 7,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ele_1273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1366_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1271_branch_req_0," req0 do_while_stmt_1271_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1271_branch_ack_0," ack0 do_while_stmt_1271_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1271_branch_ack_1," ack1 do_while_stmt_1271_branch");
    do_while_stmt_1271_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u7_u1_1399_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1271_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1271_branch_req_0,
          ack0 => do_while_stmt_1271_branch_ack_0,
          ack1 => do_while_stmt_1271_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1248_branch_req_0," req0 if_stmt_1248_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1248_branch_ack_0," ack0 if_stmt_1248_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1248_branch_ack_1," ack1 if_stmt_1248_branch");
    if_stmt_1248_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u16_u1_1251_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1248_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1248_branch_req_0,
          ack0 => if_stmt_1248_branch_ack_0,
          ack1 => if_stmt_1248_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1266_branch_req_0," req0 if_stmt_1266_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1266_branch_ack_0," ack0 if_stmt_1266_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1266_branch_ack_1," ack1 if_stmt_1266_branch");
    if_stmt_1266_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u2_u1_1269_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1266_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1266_branch_req_0,
          ack0 => if_stmt_1266_branch_ack_0,
          ack1 => if_stmt_1266_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u16_u16_1255_inst flow-through 
    process(n_iter_1256) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ADD_u16_u16_1255_inst:flowthrough inputs: " & " iter_1239 = "& Convert_SLV_To_Hex_String(iter_1239) & " konst_1254_wire_constant = "& Convert_SLV_To_Hex_String(konst_1254_wire_constant) & " outputs:" & " n_iter_1256= "  & Convert_SLV_To_Hex_String(n_iter_1256));
      --
    end process; 
    -- binary operator ADD_u16_u16_1255_inst
    process(iter_1239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iter_1239, konst_1254_wire_constant, tmp_var);
      n_iter_1256 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u5_u5_1320_inst flow-through 
    process(ADD_u5_u5_1320_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ADD_u5_u5_1320_inst:flowthrough inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " konst_1319_wire_constant = "& Convert_SLV_To_Hex_String(konst_1319_wire_constant) & " outputs:" & " ADD_u5_u5_1320_wire= "  & Convert_SLV_To_Hex_String(ADD_u5_u5_1320_wire));
      --
    end process; 
    -- binary operator ADD_u5_u5_1320_inst
    process(J_1279) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntAdd_proc(J_1279, konst_1319_wire_constant, tmp_var);
      ADD_u5_u5_1320_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_1298_inst flow-through 
    process(ADD_u6_u6_1298_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ADD_u6_u6_1298_inst:flowthrough inputs: " & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " konst_1297_wire_constant = "& Convert_SLV_To_Hex_String(konst_1297_wire_constant) & " outputs:" & " ADD_u6_u6_1298_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_1298_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_1298_inst
    process(I_1284) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_1284, konst_1297_wire_constant, tmp_var);
      ADD_u6_u6_1298_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_1331_inst flow-through 
    process(ADD_u6_u6_1331_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ADD_u6_u6_1331_inst:flowthrough inputs: " & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " konst_1330_wire_constant = "& Convert_SLV_To_Hex_String(konst_1330_wire_constant) & " outputs:" & " ADD_u6_u6_1331_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_1331_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_1331_inst
    process(I_1284) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_1284, konst_1330_wire_constant, tmp_var);
      ADD_u6_u6_1331_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u7_u7_1311_inst flow-through 
    process(ADD_u7_u7_1311_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ADD_u7_u7_1311_inst:flowthrough inputs: " & " ele_1273 = "& Convert_SLV_To_Hex_String(ele_1273) & " konst_1310_wire_constant = "& Convert_SLV_To_Hex_String(konst_1310_wire_constant) & " outputs:" & " ADD_u7_u7_1311_wire= "  & Convert_SLV_To_Hex_String(ADD_u7_u7_1311_wire));
      --
    end process; 
    -- binary operator ADD_u7_u7_1311_inst
    process(ele_1273) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ele_1273, konst_1310_wire_constant, tmp_var);
      ADD_u7_u7_1311_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u16_u1_1251_inst flow-through 
    process(EQ_u16_u1_1251_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:EQ_u16_u1_1251_inst:flowthrough inputs: " & " cmd_1247 = "& Convert_SLV_To_Hex_String(cmd_1247) & " iter_1239 = "& Convert_SLV_To_Hex_String(iter_1239) & " outputs:" & " EQ_u16_u1_1251_wire= "  & Convert_SLV_To_Hex_String(EQ_u16_u1_1251_wire));
      --
    end process; 
    -- binary operator EQ_u16_u1_1251_inst
    process(cmd_1247, iter_1239) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(cmd_1247, iter_1239, tmp_var);
      EQ_u16_u1_1251_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1269_inst flow-through 
    process(EQ_u2_u1_1269_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:EQ_u2_u1_1269_inst:flowthrough inputs: " & " check_both_1263 = "& Convert_SLV_To_Hex_String(check_both_1263) & " konst_1268_wire_constant = "& Convert_SLV_To_Hex_String(konst_1268_wire_constant) & " outputs:" & " EQ_u2_u1_1269_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1269_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1269_inst
    process(check_both_1263) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(check_both_1263, konst_1268_wire_constant, tmp_var);
      EQ_u2_u1_1269_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u5_u1_1328_inst flow-through 
    process(EQ_u5_u1_1328_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:EQ_u5_u1_1328_inst:flowthrough inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " konst_1327_wire_constant = "& Convert_SLV_To_Hex_String(konst_1327_wire_constant) & " outputs:" & " EQ_u5_u1_1328_wire= "  & Convert_SLV_To_Hex_String(EQ_u5_u1_1328_wire));
      --
    end process; 
    -- binary operator EQ_u5_u1_1328_inst
    process(J_1279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_1279, konst_1327_wire_constant, tmp_var);
      EQ_u5_u1_1328_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u6_u1_1351_inst flow-through 
    process(EQ_u6_u1_1351_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:EQ_u6_u1_1351_inst:flowthrough inputs: " & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " konst_1350_wire_constant = "& Convert_SLV_To_Hex_String(konst_1350_wire_constant) & " outputs:" & " EQ_u6_u1_1351_wire= "  & Convert_SLV_To_Hex_String(EQ_u6_u1_1351_wire));
      --
    end process; 
    -- binary operator EQ_u6_u1_1351_inst
    process(I_1284) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_1284, konst_1350_wire_constant, tmp_var);
      EQ_u6_u1_1351_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u5_u1_1317_inst flow-through 
    process(ULT_u5_u1_1317_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ULT_u5_u1_1317_inst:flowthrough inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " konst_1316_wire_constant = "& Convert_SLV_To_Hex_String(konst_1316_wire_constant) & " outputs:" & " ULT_u5_u1_1317_wire= "  & Convert_SLV_To_Hex_String(ULT_u5_u1_1317_wire));
      --
    end process; 
    -- binary operator ULT_u5_u1_1317_inst
    process(J_1279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(J_1279, konst_1316_wire_constant, tmp_var);
      ULT_u5_u1_1317_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u7_u1_1399_inst flow-through 
    process(ULT_u7_u1_1399_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:ULT_u7_u1_1399_inst:flowthrough inputs: " & " ele_1273 = "& Convert_SLV_To_Hex_String(ele_1273) & " konst_1398_wire_constant = "& Convert_SLV_To_Hex_String(konst_1398_wire_constant) & " outputs:" & " ULT_u7_u1_1399_wire= "  & Convert_SLV_To_Hex_String(ULT_u7_u1_1399_wire));
      --
    end process; 
    -- binary operator ULT_u7_u1_1399_inst
    process(ele_1273) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(ele_1273, konst_1398_wire_constant, tmp_var);
      ULT_u7_u1_1399_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_start_accelerator_1246_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_start_accelerator_1246_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:RPIPE_start_accelerator_1246_inst:started:   PipeRead from start_accelerator inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_start_accelerator_1246_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:RPIPE_start_accelerator_1246_inst:finished:  outputs: " & " cmd_1247= "  & Convert_SLV_To_Hex_String(cmd_1247));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_start_accelerator_1246_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_start_accelerator_1246_inst_req_0;
      RPIPE_start_accelerator_1246_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_start_accelerator_1246_inst_req_1;
      RPIPE_start_accelerator_1246_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_1247 <= data_out(15 downto 0);
      start_accelerator_read_0_gI: SplitGuardInterface generic map(name => "start_accelerator_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      start_accelerator_read_0: InputPortRevised -- 
        generic map ( name => "start_accelerator_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => start_accelerator_pipe_read_req(0),
          oack => start_accelerator_pipe_read_ack(0),
          odata => start_accelerator_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_accelerator_done_1401_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_accelerator_done_1401_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:WPIPE_accelerator_done_1401_inst:started:   PipeWrite to accelerator_done inputs: " & " type_cast_1403_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1403_wire_constant));
          --
        end if; 
        if WPIPE_accelerator_done_1401_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:WPIPE_accelerator_done_1401_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_accelerator_done_1401_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_accelerator_done_1401_inst_req_0;
      WPIPE_accelerator_done_1401_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_accelerator_done_1401_inst_req_1;
      WPIPE_accelerator_done_1401_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1403_wire_constant;
      accelerator_done_write_0_gI: SplitGuardInterface generic map(name => "accelerator_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      accelerator_done_write_0: OutputPortRevised -- 
        generic map ( name => "accelerator_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => accelerator_done_pipe_write_req(0),
          oack => accelerator_done_pipe_write_ack(0),
          odata => accelerator_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_read_sums_1364_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_read_sums_1364_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:WPIPE_read_sums_1364_inst:started:   PipeWrite to read_sums inputs: " & " type_cast_1366_wire = "& Convert_SLV_To_Hex_String(type_cast_1366_wire));
          --
        end if; 
        if WPIPE_read_sums_1364_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:WPIPE_read_sums_1364_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_read_sums_1364_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_read_sums_1364_inst_req_0;
      WPIPE_read_sums_1364_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_read_sums_1364_inst_req_1;
      WPIPE_read_sums_1364_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1366_wire;
      read_sums_write_1_gI: SplitGuardInterface generic map(name => "read_sums_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      read_sums_write_1: OutputPortRevised -- 
        generic map ( name => "read_sums", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => read_sums_pipe_write_req(0),
          oack => read_sums_pipe_write_ack(0),
          odata => read_sums_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator call_stmt_1259_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1259_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1259_call:started:  Call to module initFilter inputs: " & " R_filter_start_addr_1257_wire_constant = "& Convert_SLV_To_Hex_String(R_filter_start_addr_1257_wire_constant));
          --
        end if; 
        if call_stmt_1259_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1259_call:finished:  outputs: " & " initialized_filter_1259= "  & Convert_SLV_To_Hex_String(initialized_filter_1259));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1259_call 
    initFilter_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1259_call_req_0;
      call_stmt_1259_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1259_call_req_1;
      call_stmt_1259_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initFilter_call_group_0_gI: SplitGuardInterface generic map(name => "initFilter_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_filter_start_addr_1257_wire_constant;
      initialized_filter_1259 <= data_out(1 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => initFilter_call_reqs(0),
          ackR => initFilter_call_acks(0),
          dataR => initFilter_call_data(5 downto 0),
          tagR => initFilter_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 2,
          owidth => 2,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => initFilter_return_acks(0), -- cross-over
          ackL => initFilter_return_reqs(0), -- cross-over
          dataL => initFilter_return_data(1 downto 0),
          tagL => initFilter_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1307_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1307_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1307_call:started:  Call to module initIfMaps inputs: " & " type_cast_1302_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1302_wire_constant) & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " col_to_be_replaced_1289 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1289));
          --
        end if; 
        if call_stmt_1307_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1307_call:finished:  outputs: " & " initialized_ifmaps_1307= "  & Convert_SLV_To_Hex_String(initialized_ifmaps_1307));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1307_call 
    initIfMaps_call_group_1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1307_call_req_0;
      call_stmt_1307_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1307_call_req_1;
      call_stmt_1307_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      initIfMaps_call_group_1_gI: SplitGuardInterface generic map(name => "initIfMaps_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1302_wire_constant & I_1284 & J_1279 & col_to_be_replaced_1289;
      initialized_ifmaps_1307 <= data_out(1 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 14,
        owidth => 14,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => initIfMaps_call_reqs(0),
          ackR => initIfMaps_call_acks(0),
          dataR => initIfMaps_call_data(13 downto 0),
          tagR => initIfMaps_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 2,
          owidth => 2,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => initIfMaps_return_acks(0), -- cross-over
          ackL => initIfMaps_return_reqs(0), -- cross-over
          dataL => initIfMaps_return_data(1 downto 0),
          tagL => initIfMaps_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_1339_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1339_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1339_call:started:  Call to module cal_col_to_be_replaced inputs: " & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " col_to_be_replaced_1289 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1289));
          --
        end if; 
        if call_stmt_1339_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1339_call:finished:  outputs: " & " new_col_to_be_replaced_1339= "  & Convert_SLV_To_Hex_String(new_col_to_be_replaced_1339));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_1339_call 
    cal_col_to_be_replaced_call_group_2: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1339_call_req_0;
      call_stmt_1339_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1339_call_req_1;
      call_stmt_1339_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      cal_col_to_be_replaced_call_group_2_gI: SplitGuardInterface generic map(name => "cal_col_to_be_replaced_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= J_1279 & col_to_be_replaced_1289;
      new_col_to_be_replaced_1339 <= data_out(1 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 7,
        owidth => 7,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => cal_col_to_be_replaced_call_reqs(0),
          ackR => cal_col_to_be_replaced_call_acks(0),
          dataR => cal_col_to_be_replaced_call_data(6 downto 0),
          tagR => cal_col_to_be_replaced_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 2,
          owidth => 2,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => cal_col_to_be_replaced_return_acks(0), -- cross-over
          ackL => cal_col_to_be_replaced_return_reqs(0), -- cross-over
          dataL => cal_col_to_be_replaced_return_data(1 downto 0),
          tagL => cal_col_to_be_replaced_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_1347_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1347_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1347_call:started:  Call to module mainAcc inputs: " & " I_1284 = "& Convert_SLV_To_Hex_String(I_1284) & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " col_to_be_replaced_1289 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1289));
          --
        end if; 
        if call_stmt_1347_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1347_call:finished:  outputs: " & " ofmap_pixel_1347= "  & Convert_SLV_To_Hex_String(ofmap_pixel_1347));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_1347_call 
    mainAcc_call_group_3: Block -- 
      signal data_in: std_logic_vector(12 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1347_call_req_0;
      call_stmt_1347_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1347_call_req_1;
      call_stmt_1347_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      mainAcc_call_group_3_gI: SplitGuardInterface generic map(name => "mainAcc_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= I_1284 & J_1279 & col_to_be_replaced_1289;
      ofmap_pixel_1347 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 13,
        owidth => 13,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => mainAcc_call_reqs(0),
          ackR => mainAcc_call_acks(0),
          dataR => mainAcc_call_data(12 downto 0),
          tagR => mainAcc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => mainAcc_return_acks(0), -- cross-over
          ackL => mainAcc_return_reqs(0), -- cross-over
          dataL => mainAcc_return_data(15 downto 0),
          tagL => mainAcc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- logger for split-operator call_stmt_1363_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1363_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1363_call:started:  Call to module mainAcc2 inputs: " & " checkIFour_1357 (guard complement )= " & Convert_SLV_To_String(checkIFour_1357) & " I_1_1300 = "& Convert_SLV_To_Hex_String(I_1_1300) & " J_1279 = "& Convert_SLV_To_Hex_String(J_1279) & " col_to_be_replaced_1289 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1289));
          --
        end if; 
        if call_stmt_1363_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1363_call:finished:  outputs: " & " ofmap_pixel2_1363= "  & Convert_SLV_To_Hex_String(ofmap_pixel2_1363));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (4) : call_stmt_1363_call 
    mainAcc2_call_group_4: Block -- 
      signal data_in: std_logic_vector(12 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1363_call_req_0;
      call_stmt_1363_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1363_call_req_1;
      call_stmt_1363_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not checkIFour_1357(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      mainAcc2_call_group_4_gI: SplitGuardInterface generic map(name => "mainAcc2_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= I_1_1300 & J_1279 & col_to_be_replaced_1289;
      ofmap_pixel2_1363 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 13,
        owidth => 13,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => mainAcc2_call_reqs(0),
          ackR => mainAcc2_call_acks(0),
          dataR => mainAcc2_call_data(12 downto 0),
          tagR => mainAcc2_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => mainAcc2_return_acks(0), -- cross-over
          ackL => mainAcc2_return_reqs(0), -- cross-over
          dataL => mainAcc2_return_data(15 downto 0),
          tagL => mainAcc2_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- logger for split-operator call_stmt_1379_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1379_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1379_call:started:  Call to module accessMem inputs: " & " R_write_signal_1374_wire_constant = "& Convert_SLV_To_Hex_String(R_write_signal_1374_wire_constant) & " I_1457_delayed_4_0_1370 = "& Convert_SLV_To_Hex_String(I_1457_delayed_4_0_1370) & " J_1458_delayed_4_0_1373 = "& Convert_SLV_To_Hex_String(J_1458_delayed_4_0_1373) & " ofmap_pixel_1347 = "& Convert_SLV_To_Hex_String(ofmap_pixel_1347));
          --
        end if; 
        if call_stmt_1379_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1379_call:finished:  outputs: " & " r_data_sum_cal_1379= "  & Convert_SLV_To_Hex_String(r_data_sum_cal_1379));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_1395_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1395_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1395_call:started:  Call to module accessMem inputs: " & " checkIFour_1462_delayed_4_0_1382 (guard complement )= " & Convert_SLV_To_String(checkIFour_1462_delayed_4_0_1382) & " R_write_signal_1390_wire_constant = "& Convert_SLV_To_Hex_String(R_write_signal_1390_wire_constant) & " I_1_1464_delayed_4_0_1385 = "& Convert_SLV_To_Hex_String(I_1_1464_delayed_4_0_1385) & " J_1465_delayed_4_0_1388 = "& Convert_SLV_To_Hex_String(J_1465_delayed_4_0_1388) & " ofmap_pixel2_1363 = "& Convert_SLV_To_Hex_String(ofmap_pixel2_1363));
          --
        end if; 
        if call_stmt_1395_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accelerator:DP:call_stmt_1395_call:finished:  outputs: " & " r_data_sum_cal2_1395= "  & Convert_SLV_To_Hex_String(r_data_sum_cal2_1395));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (5) : call_stmt_1379_call call_stmt_1395_call 
    accessMem_call_group_5: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 7, 1 => 7);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1379_call_req_0;
      reqL_unguarded(0) <= call_stmt_1395_call_req_0;
      call_stmt_1379_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1395_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1379_call_req_1;
      reqR_unguarded(0) <= call_stmt_1395_call_req_1;
      call_stmt_1379_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1395_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not checkIFour_1462_delayed_4_0_1382(0);
      guard_vector(1)  <=  '1';
      accessMem_call_group_5_accessRegulator_0: access_regulator_base generic map (name => "accessMem_call_group_5_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMem_call_group_5_accessRegulator_1: access_regulator_base generic map (name => "accessMem_call_group_5_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMem_call_group_5_gI: SplitGuardInterface generic map(name => "accessMem_call_group_5_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_write_signal_1374_wire_constant & I_1457_delayed_4_0_1370 & J_1458_delayed_4_0_1373 & ofmap_pixel_1347 & R_write_signal_1390_wire_constant & I_1_1464_delayed_4_0_1385 & J_1465_delayed_4_0_1388 & ofmap_pixel2_1363;
      r_data_sum_cal_1379 <= data_out(31 downto 16);
      r_data_sum_cal2_1395 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 56,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 5,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- 
  end Block; -- data_path
  -- 
end accelerator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    read_write_bar_1 : in  std_logic_vector(0 downto 0);
    row_index : in  std_logic_vector(5 downto 0);
    col_index : in  std_logic_vector(4 downto 0);
    write_data_1 : in  std_logic_vector(15 downto 0);
    read_data_1 : out  std_logic_vector(15 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMem;
architecture accessMem_arch of accessMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 28)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal read_write_bar_1_buffer :  std_logic_vector(0 downto 0);
  signal read_write_bar_1_update_enable: Boolean;
  signal row_index_buffer :  std_logic_vector(5 downto 0);
  signal row_index_update_enable: Boolean;
  signal col_index_buffer :  std_logic_vector(4 downto 0);
  signal col_index_update_enable: Boolean;
  signal write_data_1_buffer :  std_logic_vector(15 downto 0);
  signal write_data_1_update_enable: Boolean;
  -- output port buffer signals
  signal read_data_1_buffer :  std_logic_vector(15 downto 0);
  signal read_data_1_update_enable: Boolean;
  signal accessMem_CP_0_start: Boolean;
  signal accessMem_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_62_index_0_scale_req_0 : boolean;
  signal array_obj_ref_62_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_62_index_0_scale_req_1 : boolean;
  signal array_obj_ref_62_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_62_index_sum_1_req_0 : boolean;
  signal array_obj_ref_62_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_62_index_sum_1_req_1 : boolean;
  signal array_obj_ref_62_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_62_load_0_req_0 : boolean;
  signal array_obj_ref_62_load_0_ack_0 : boolean;
  signal array_obj_ref_62_load_0_req_1 : boolean;
  signal array_obj_ref_62_load_0_ack_1 : boolean;
  signal array_obj_ref_67_index_0_scale_req_0 : boolean;
  signal array_obj_ref_67_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_67_index_0_scale_req_1 : boolean;
  signal array_obj_ref_67_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_67_index_sum_1_req_0 : boolean;
  signal array_obj_ref_67_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_67_index_sum_1_req_1 : boolean;
  signal array_obj_ref_67_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_67_store_0_req_0 : boolean;
  signal array_obj_ref_67_store_0_ack_0 : boolean;
  signal array_obj_ref_67_store_0_req_1 : boolean;
  signal array_obj_ref_67_store_0_ack_1 : boolean;
  signal W_read_write_bar_1_71_delayed_4_0_70_inst_req_0 : boolean;
  signal W_read_write_bar_1_71_delayed_4_0_70_inst_ack_0 : boolean;
  signal W_read_write_bar_1_71_delayed_4_0_70_inst_req_1 : boolean;
  signal W_read_write_bar_1_71_delayed_4_0_70_inst_ack_1 : boolean;
  signal MUX_77_inst_req_0 : boolean;
  signal MUX_77_inst_ack_0 : boolean;
  signal MUX_77_inst_req_1 : boolean;
  signal MUX_77_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMem_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 28) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= read_write_bar_1;
  read_write_bar_1_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(6 downto 1) <= row_index;
  row_index_buffer <= in_buffer_data_out(6 downto 1);
  in_buffer_data_in(11 downto 7) <= col_index;
  col_index_buffer <= in_buffer_data_out(11 downto 7);
  in_buffer_data_in(27 downto 12) <= write_data_1;
  write_data_1_buffer <= in_buffer_data_out(27 downto 12);
  in_buffer_data_in(tag_length + 27 downto 28) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 27 downto 28);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 5) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 1,5 => 7);
    constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 7);
    constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 6); -- 
  begin -- 
    preds <= read_write_bar_1_update_enable & row_index_update_enable & col_index_update_enable & write_data_1_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMem_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= read_data_1_buffer;
  read_data_1 <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  read_data_1_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "read_data_1_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_read_data_1_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => read_data_1_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMem_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_start,"accessMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMem_CP_0_symbol, "accessMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMem_CP_0: Block -- control-path 
    signal accessMem_CP_0_elements: BooleanArray(48 downto 0);
    -- 
  begin -- 
    accessMem_CP_0_elements(0) <= accessMem_CP_0_start;
    accessMem_CP_0_symbol <= accessMem_CP_0_elements(48);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessMem_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	15 
    -- CP-element group 1: 	20 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	27 
    -- CP-element group 1: 	28 
    -- CP-element group 1: 	33 
    -- CP-element group 1:  members (35) 
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resized_0
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_computed_0
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resized_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_computed_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resized_0
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_computed_0
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resized_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_computed_1
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_1/scale_rename_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(1) <= accessMem_CP_0_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	35 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	43 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_63_to_assign_stmt_78/read_write_bar_1_update_enable
      -- CP-element group 2: 	 assign_stmt_63_to_assign_stmt_78/read_write_bar_1_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(18) & accessMem_CP_0_elements(31) & accessMem_CP_0_elements(35);
      gj_accessMem_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: 	22 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_63_to_assign_stmt_78/row_index_update_enable
      -- CP-element group 3: 	 assign_stmt_63_to_assign_stmt_78/row_index_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(9) & accessMem_CP_0_elements(22);
      gj_accessMem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	29 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	45 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_63_to_assign_stmt_78/col_index_update_enable
      -- CP-element group 4: 	 assign_stmt_63_to_assign_stmt_78/col_index_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(16) & accessMem_CP_0_elements(29);
      gj_accessMem_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	31 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	46 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_63_to_assign_stmt_78/write_data_1_update_enable
      -- CP-element group 5: 	 assign_stmt_63_to_assign_stmt_78/write_data_1_update_enable_out
      -- 
    -- logger for CP element group accessMem_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(31);
      gj_accessMem_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	47 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	38 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_63_to_assign_stmt_78/read_data_1_update_enable
      -- CP-element group 6: 	 assign_stmt_63_to_assign_stmt_78/read_data_1_update_enable_in
      -- 
    -- logger for CP element group accessMem_CP_0_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(6) <= accessMem_CP_0_elements(47);
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: 	17 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	18 
    -- CP-element group 7: 	31 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	18 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_sample_start_
      -- CP-element group 7: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/$entry
      -- CP-element group 7: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/$entry
      -- CP-element group 7: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_97_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_97_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(7), ack => array_obj_ref_62_load_0_req_0); -- 
    accessMem_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(17) & accessMem_CP_0_elements(18) & accessMem_CP_0_elements(31);
      gj_accessMem_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	19 
    -- CP-element group 8: 	39 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_update_start_
      -- CP-element group 8: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/$entry
      -- CP-element group 8: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/$entry
      -- CP-element group 8: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/word_0/$entry
      -- CP-element group 8: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(8), ack => array_obj_ref_62_load_0_req_1); -- 
    accessMem_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(19) & accessMem_CP_0_elements(39);
      gj_accessMem_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	3 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scaled_0
      -- 
    -- logger for CP element group accessMem_CP_0_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "accessMem_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(13) & accessMem_CP_0_elements(16);
      gj_accessMem_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_sample_start
      -- CP-element group 10: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_0_scale_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_39_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_39_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(10), ack => array_obj_ref_62_index_0_scale_req_0); -- 
    accessMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(12);
      gj_accessMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_update_start
      -- CP-element group 11: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Update/$entry
      -- CP-element group 11: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_0_scale_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(11), ack => array_obj_ref_62_index_0_scale_req_1); -- 
    accessMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(13);
      gj_accessMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	42 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_sample_complete
      -- CP-element group 12: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_0_scale_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_40_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_0_scale_ack_0, ack => accessMem_CP_0_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_update_complete
      -- CP-element group 13: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Update/$exit
      -- CP-element group 13: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_index_scale_0_Update/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_0_scale_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_45_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_0_scale_ack_1, ack => accessMem_CP_0_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_sample_start
      -- CP-element group 14: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_sum_1_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(14), ack => array_obj_ref_62_index_sum_1_req_0); -- 
    accessMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(9) & accessMem_CP_0_elements(16);
      gj_accessMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_update_start
      -- CP-element group 15: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Update/$entry
      -- CP-element group 15: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_sum_1_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(15), ack => array_obj_ref_62_index_sum_1_req_1); -- 
    accessMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(17) & accessMem_CP_0_elements(18);
      gj_accessMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	42 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_sample_complete
      -- CP-element group 16: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_sum_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_sum_1_ack_0, ack => accessMem_CP_0_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	7 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (18) 
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_word_address_calculated
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_root_address_calculated
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_offset_calculated
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_update_complete
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Update/$exit
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_partial_sum_1_Update/ca
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_final_index_sum_regn/$entry
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_final_index_sum_regn/$exit
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_final_index_sum_regn/req
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_final_index_sum_regn/ack
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_base_plus_offset/$entry
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_base_plus_offset/$exit
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_word_addrgen/$entry
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_word_addrgen/$exit
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_word_addrgen/root_register_req
      -- CP-element group 17: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_index_sum_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_sum_1_ack_1, ack => accessMem_CP_0_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	7 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: 	7 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_sample_completed_
      -- CP-element group 18: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/$exit
      -- CP-element group 18: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/word_0/$exit
      -- CP-element group 18: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_98_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_load_0_ack_0, ack => accessMem_CP_0_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	37 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	8 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_update_completed_
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/$exit
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/$exit
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/word_0/$exit
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/word_access_complete/word_0/ca
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/array_obj_ref_62_Merge/$entry
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/array_obj_ref_62_Merge/$exit
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/array_obj_ref_62_Merge/merge_req
      -- CP-element group 19: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_Update/array_obj_ref_62_Merge/merge_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_62_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_load_0_ack_1, ack => accessMem_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: 	30 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	31 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_sample_start_
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/$entry
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/array_obj_ref_67_Split/$entry
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/array_obj_ref_67_Split/$exit
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/array_obj_ref_67_Split/split_req
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/array_obj_ref_67_Split/split_ack
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/$entry
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(20), ack => array_obj_ref_67_store_0_req_0); -- 
    accessMem_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(30) & accessMem_CP_0_elements(41) & accessMem_CP_0_elements(31);
      gj_accessMem_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	32 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_update_start_
      -- CP-element group 21: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/$entry
      -- CP-element group 21: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/$entry
      -- CP-element group 21: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/word_0/$entry
      -- CP-element group 21: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(21), ack => array_obj_ref_67_store_0_req_1); -- 
    accessMem_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMem_CP_0_elements(32);
      gj_accessMem_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	29 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	3 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scaled_0
      -- 
    -- logger for CP element group accessMem_CP_0_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(26) & accessMem_CP_0_elements(29);
      gj_accessMem_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_sample_start
      -- CP-element group 23: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_0_scale_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(23), ack => array_obj_ref_67_index_0_scale_req_0); -- 
    accessMem_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(25);
      gj_accessMem_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_update_start
      -- CP-element group 24: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Update/$entry
      -- CP-element group 24: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_0_scale_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(24), ack => array_obj_ref_67_index_0_scale_req_1); -- 
    accessMem_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(26);
      gj_accessMem_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	42 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_sample_complete
      -- CP-element group 25: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_0_scale_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_0_scale_ack_0, ack => accessMem_CP_0_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_update_complete
      -- CP-element group 26: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Update/$exit
      -- CP-element group 26: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_index_scale_0_Update/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_0_scale_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_0_scale_ack_1, ack => accessMem_CP_0_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: 	22 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_sample_start
      -- CP-element group 27: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Sample/rr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_sum_1_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(27), ack => array_obj_ref_67_index_sum_1_req_0); -- 
    accessMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(22) & accessMem_CP_0_elements(29);
      gj_accessMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	1 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: 	31 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_update_start
      -- CP-element group 28: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Update/$entry
      -- CP-element group 28: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Update/cr
      -- 
    -- logger for CP element group accessMem_CP_0_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_sum_1_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(28), ack => array_obj_ref_67_index_sum_1_req_1); -- 
    accessMem_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(30) & accessMem_CP_0_elements(31);
      gj_accessMem_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	42 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_sample_complete
      -- CP-element group 29: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Sample/ra
      -- 
    -- logger for CP element group accessMem_CP_0_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_sum_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_sum_1_ack_0, ack => accessMem_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	20 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (18) 
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_word_address_calculated
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_root_address_calculated
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_offset_calculated
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_update_complete
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Update/$exit
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_partial_sum_1_Update/ca
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_final_index_sum_regn/$entry
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_final_index_sum_regn/$exit
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_final_index_sum_regn/req
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_final_index_sum_regn/ack
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_base_plus_offset/$entry
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_base_plus_offset/$exit
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_word_addrgen/$entry
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_word_addrgen/$exit
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_word_addrgen/root_register_req
      -- CP-element group 30: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_index_sum_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_index_sum_1_ack_1, ack => accessMem_CP_0_elements(30)); -- 
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	20 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	42 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: 	5 
    -- CP-element group 31: 	7 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	28 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_sample_completed_
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/$exit
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Sample/word_access_start/word_0/ra
      -- CP-element group 31: 	 assign_stmt_63_to_assign_stmt_78/ring_reenable_memory_space_3
      -- 
    -- logger for CP element group accessMem_CP_0_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_store_0_ack_0, ack => accessMem_CP_0_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	21 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	42 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	21 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_update_completed_
      -- CP-element group 32: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/$exit
      -- CP-element group 32: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/$exit
      -- CP-element group 32: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_67_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group accessMem_CP_0_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:array_obj_ref_67_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_67_store_0_ack_1, ack => accessMem_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	1 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_sample_start_
      -- CP-element group 33: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Sample/$entry
      -- CP-element group 33: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Sample/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_1_71_delayed_4_0_70_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(33), ack => W_read_write_bar_1_71_delayed_4_0_70_inst_req_0); -- 
    accessMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(1) & accessMem_CP_0_elements(35);
      gj_accessMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	39 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_update_start_
      -- CP-element group 34: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Update/$entry
      -- CP-element group 34: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Update/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_1_71_delayed_4_0_70_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(34), ack => W_read_write_bar_1_71_delayed_4_0_70_inst_req_1); -- 
    accessMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(36) & accessMem_CP_0_elements(39);
      gj_accessMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	2 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_sample_completed_
      -- CP-element group 35: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Sample/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_1_71_delayed_4_0_70_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_1_71_delayed_4_0_70_inst_ack_0, ack => accessMem_CP_0_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_update_completed_
      -- CP-element group 36: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Update/$exit
      -- CP-element group 36: 	 assign_stmt_63_to_assign_stmt_78/assign_stmt_72_Update/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:W_read_write_bar_1_71_delayed_4_0_70_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_write_bar_1_71_delayed_4_0_70_inst_ack_1, ack => accessMem_CP_0_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	19 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_sample_start_
      -- CP-element group 37: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_start/$entry
      -- CP-element group 37: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_start/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_77_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(37), ack => MUX_77_inst_req_0); -- 
    accessMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(19) & accessMem_CP_0_elements(36) & accessMem_CP_0_elements(39);
      gj_accessMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	6 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_update_start_
      -- CP-element group 38: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_complete/$entry
      -- CP-element group 38: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_complete/req
      -- 
    -- logger for CP element group accessMem_CP_0_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_77_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMem_CP_0_elements(38), ack => MUX_77_inst_req_1); -- 
    accessMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(6) & accessMem_CP_0_elements(40);
      gj_accessMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	8 
    -- CP-element group 39: 	34 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_sample_completed_
      -- CP-element group 39: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_start/$exit
      -- CP-element group 39: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_start/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_77_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_77_inst_ack_0, ack => accessMem_CP_0_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_update_completed_
      -- CP-element group 40: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_complete/$exit
      -- CP-element group 40: 	 assign_stmt_63_to_assign_stmt_78/MUX_77_complete/ack
      -- 
    -- logger for CP element group accessMem_CP_0_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:MUX_77_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_77_inst_ack_1, ack => accessMem_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 assign_stmt_63_to_assign_stmt_78/array_obj_ref_62_array_obj_ref_67_delay
      -- 
    -- logger for CP element group accessMem_CP_0_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group accessMem_CP_0_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => accessMem_CP_0_elements(18), ack => accessMem_CP_0_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	12 
    -- CP-element group 42: 	16 
    -- CP-element group 42: 	25 
    -- CP-element group 42: 	29 
    -- CP-element group 42: 	31 
    -- CP-element group 42: 	32 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	48 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 assign_stmt_63_to_assign_stmt_78/$exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "accessMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= accessMem_CP_0_elements(12) & accessMem_CP_0_elements(16) & accessMem_CP_0_elements(25) & accessMem_CP_0_elements(29) & accessMem_CP_0_elements(31) & accessMem_CP_0_elements(32) & accessMem_CP_0_elements(40);
      gj_accessMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMem_CP_0_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  place  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	2 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 read_write_bar_1_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(43) <= accessMem_CP_0_elements(2);
    -- CP-element group 44:  place  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 row_index_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(44) <= accessMem_CP_0_elements(3);
    -- CP-element group 45:  place  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	4 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 col_index_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(45) <= accessMem_CP_0_elements(4);
    -- CP-element group 46:  place  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	5 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 write_data_1_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(46) <= accessMem_CP_0_elements(5);
    -- CP-element group 47:  place  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	6 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 read_data_1_update_enable
      -- 
    -- logger for CP element group accessMem_CP_0_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 48:  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	42 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 $exit
      -- 
    -- logger for CP element group accessMem_CP_0_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMem_CP_0_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMem:CP:accessMem_CP_0_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    accessMem_CP_0_elements(48) <= accessMem_CP_0_elements(42);
    --  hookup: inputs to control-path 
    accessMem_CP_0_elements(47) <= read_data_1_update_enable;
    -- hookup: output from control-path 
    read_write_bar_1_update_enable <= accessMem_CP_0_elements(43);
    row_index_update_enable <= accessMem_CP_0_elements(44);
    col_index_update_enable <= accessMem_CP_0_elements(45);
    write_data_1_update_enable <= accessMem_CP_0_elements(46);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_col_index_61_resized : std_logic_vector(6 downto 0);
    signal R_col_index_61_scaled : std_logic_vector(6 downto 0);
    signal R_col_index_66_resized : std_logic_vector(6 downto 0);
    signal R_col_index_66_scaled : std_logic_vector(6 downto 0);
    signal R_row_index_60_resized : std_logic_vector(6 downto 0);
    signal R_row_index_60_scaled : std_logic_vector(6 downto 0);
    signal R_row_index_65_resized : std_logic_vector(6 downto 0);
    signal R_row_index_65_scaled : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_62_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_index_partial_sum_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_word_address_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_62_word_offset_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_67_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_index_partial_sum_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_word_address_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_67_word_offset_0 : std_logic_vector(6 downto 0);
    signal konst_76_wire_constant : std_logic_vector(15 downto 0);
    signal read_write_bar_1_71_delayed_4_0_72 : std_logic_vector(0 downto 0);
    signal t_read_data_11_63 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_62_offset_scale_factor_0 <= "0001000";
    array_obj_ref_62_offset_scale_factor_1 <= "0000001";
    array_obj_ref_62_resized_base_address <= "0000000";
    array_obj_ref_62_word_offset_0 <= "0000000";
    array_obj_ref_67_offset_scale_factor_0 <= "0001000";
    array_obj_ref_67_offset_scale_factor_1 <= "0000001";
    array_obj_ref_67_resized_base_address <= "0000000";
    array_obj_ref_67_word_offset_0 <= "0000000";
    konst_76_wire_constant <= "0000000000000000";
    -- logger for split-operator MUX_77_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_77_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_77_inst:started:   inputs: " & " read_write_bar_1_71_delayed_4_0_72 = "& Convert_SLV_To_Hex_String(read_write_bar_1_71_delayed_4_0_72) & " t_read_data_11_63 = "& Convert_SLV_To_Hex_String(t_read_data_11_63) & " konst_76_wire_constant = "& Convert_SLV_To_Hex_String(konst_76_wire_constant));
          --
        end if; 
        if MUX_77_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:MUX_77_inst:finished:  outputs: " & " read_data_1_buffer= "  & Convert_SLV_To_Hex_String(read_data_1_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_77_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_77_inst_req_0;
      MUX_77_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_77_inst_req_1;
      MUX_77_inst_ack_1<= update_ack(0);
      MUX_77_inst: SelectSplitProtocol generic map(name => "MUX_77_inst", data_width => 16, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => t_read_data_11_63, y => konst_76_wire_constant, sel => read_write_bar_1_71_delayed_4_0_72, z => read_data_1_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator W_read_write_bar_1_71_delayed_4_0_70_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_read_write_bar_1_71_delayed_4_0_70_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_1_71_delayed_4_0_70_inst:started:   inputs: " & " read_write_bar_1_buffer = "& Convert_SLV_To_Hex_String(read_write_bar_1_buffer));
          --
        end if; 
        if W_read_write_bar_1_71_delayed_4_0_70_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:W_read_write_bar_1_71_delayed_4_0_70_inst:finished:  outputs: " & " read_write_bar_1_71_delayed_4_0_72= "  & Convert_SLV_To_Hex_String(read_write_bar_1_71_delayed_4_0_72));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_read_write_bar_1_71_delayed_4_0_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_write_bar_1_71_delayed_4_0_70_inst_req_0;
      W_read_write_bar_1_71_delayed_4_0_70_inst_ack_0<= wack(0);
      rreq(0) <= W_read_write_bar_1_71_delayed_4_0_70_inst_req_1;
      W_read_write_bar_1_71_delayed_4_0_70_inst_ack_1<= rack(0);
      W_read_write_bar_1_71_delayed_4_0_70_inst : InterlockBuffer generic map ( -- 
        name => "W_read_write_bar_1_71_delayed_4_0_70_inst",
        buffer_size => 4,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_write_bar_1_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_write_bar_1_71_delayed_4_0_72,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_62_addr_0 flow-through 
    process(array_obj_ref_62_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_addr_0:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_62_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_62_root_address) & "outputs: " & " array_obj_ref_62_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_62_addr_0
    process(array_obj_ref_62_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_root_address;
      ov(6 downto 0) := iv;
      array_obj_ref_62_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_gather_scatter flow-through 
    process(t_read_data_11_63) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_gather_scatter:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_62_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_62_data_0) & "outputs: " & " t_read_data_11_63= "  & Convert_SLV_To_Hex_String(t_read_data_11_63));
      --
    end process; 
    -- equivalence array_obj_ref_62_gather_scatter
    process(array_obj_ref_62_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_data_0;
      ov(15 downto 0) := iv;
      t_read_data_11_63 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_index_0_resize flow-through 
    process(R_row_index_60_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_0_resize:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " row_index_buffer = "& Convert_SLV_To_Hex_String(row_index_buffer) & "outputs: " & " R_row_index_60_resized= "  & Convert_SLV_To_Hex_String(R_row_index_60_resized));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_0_resize
    process(row_index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := row_index_buffer;
      ov(5 downto 0) := iv;
      R_row_index_60_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_index_1_rename flow-through 
    process(R_col_index_61_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_1_rename:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_col_index_61_resized = "& Convert_SLV_To_Hex_String(R_col_index_61_resized) & "outputs: " & " R_col_index_61_scaled= "  & Convert_SLV_To_Hex_String(R_col_index_61_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_1_rename
    process(R_col_index_61_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_index_61_resized;
      ov(6 downto 0) := iv;
      R_col_index_61_scaled <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_index_1_resize flow-through 
    process(R_col_index_61_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_1_resize:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " col_index_buffer = "& Convert_SLV_To_Hex_String(col_index_buffer) & "outputs: " & " R_col_index_61_resized= "  & Convert_SLV_To_Hex_String(R_col_index_61_resized));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_1_resize
    process(col_index_buffer) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_index_buffer;
      ov(4 downto 0) := iv;
      R_col_index_61_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_index_offset flow-through 
    process(array_obj_ref_62_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_offset:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_62_index_partial_sum_1 = "& Convert_SLV_To_Hex_String(array_obj_ref_62_index_partial_sum_1) & "outputs: " & " array_obj_ref_62_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_62_index_offset
    process(array_obj_ref_62_index_partial_sum_1) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_index_partial_sum_1;
      ov(6 downto 0) := iv;
      array_obj_ref_62_final_offset <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_62_root_address_inst flow-through 
    process(array_obj_ref_62_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_root_address_inst:flowthrough  inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_62_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_62_final_offset) & "outputs: " & " array_obj_ref_62_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_62_root_address_inst
    process(array_obj_ref_62_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_62_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_addr_0 flow-through 
    process(array_obj_ref_67_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_addr_0:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_67_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_67_root_address) & "outputs: " & " array_obj_ref_67_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_67_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_67_addr_0
    process(array_obj_ref_67_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_67_root_address;
      ov(6 downto 0) := iv;
      array_obj_ref_67_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_gather_scatter flow-through 
    process(array_obj_ref_67_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_gather_scatter:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " write_data_1_buffer = "& Convert_SLV_To_Hex_String(write_data_1_buffer) & "outputs: " & " array_obj_ref_67_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_67_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_67_gather_scatter
    process(write_data_1_buffer) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := write_data_1_buffer;
      ov(15 downto 0) := iv;
      array_obj_ref_67_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_index_0_resize flow-through 
    process(R_row_index_65_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_0_resize:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " row_index_buffer = "& Convert_SLV_To_Hex_String(row_index_buffer) & "outputs: " & " R_row_index_65_resized= "  & Convert_SLV_To_Hex_String(R_row_index_65_resized));
      --
    end process; 
    -- equivalence array_obj_ref_67_index_0_resize
    process(row_index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := row_index_buffer;
      ov(5 downto 0) := iv;
      R_row_index_65_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_index_1_rename flow-through 
    process(R_col_index_66_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_1_rename:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_col_index_66_resized = "& Convert_SLV_To_Hex_String(R_col_index_66_resized) & "outputs: " & " R_col_index_66_scaled= "  & Convert_SLV_To_Hex_String(R_col_index_66_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_67_index_1_rename
    process(R_col_index_66_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_index_66_resized;
      ov(6 downto 0) := iv;
      R_col_index_66_scaled <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_index_1_resize flow-through 
    process(R_col_index_66_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_1_resize:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " col_index_buffer = "& Convert_SLV_To_Hex_String(col_index_buffer) & "outputs: " & " R_col_index_66_resized= "  & Convert_SLV_To_Hex_String(R_col_index_66_resized));
      --
    end process; 
    -- equivalence array_obj_ref_67_index_1_resize
    process(col_index_buffer) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_index_buffer;
      ov(4 downto 0) := iv;
      R_col_index_66_resized <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_index_offset flow-through 
    process(array_obj_ref_67_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_offset:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_67_index_partial_sum_1 = "& Convert_SLV_To_Hex_String(array_obj_ref_67_index_partial_sum_1) & "outputs: " & " array_obj_ref_67_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_67_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_67_index_offset
    process(array_obj_ref_67_index_partial_sum_1) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_67_index_partial_sum_1;
      ov(6 downto 0) := iv;
      array_obj_ref_67_final_offset <= ov(6 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_67_root_address_inst flow-through 
    process(array_obj_ref_67_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_root_address_inst:flowthrough  inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_67_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_67_final_offset) & "outputs: " & " array_obj_ref_67_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_67_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_67_root_address_inst
    process(array_obj_ref_67_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_67_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_67_root_address <= ov(6 downto 0);
      --
    end process;
    -- logger for split-operator array_obj_ref_62_index_0_scale
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_62_index_0_scale_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_0_scale:started:   inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_row_index_60_resized = "& Convert_SLV_To_Hex_String(R_row_index_60_resized) & " array_obj_ref_62_offset_scale_factor_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_62_offset_scale_factor_0));
          --
        end if; 
        if array_obj_ref_62_index_0_scale_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_0_scale:finished:  outputs: " & " R_row_index_60_scaled= "  & Convert_SLV_To_Hex_String(R_row_index_60_scaled));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_67_index_0_scale
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_67_index_0_scale_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_0_scale:started:   inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_row_index_65_resized = "& Convert_SLV_To_Hex_String(R_row_index_65_resized) & " array_obj_ref_67_offset_scale_factor_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_67_offset_scale_factor_0));
          --
        end if; 
        if array_obj_ref_67_index_0_scale_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_0_scale:finished:  outputs: " & " R_row_index_65_scaled= "  & Convert_SLV_To_Hex_String(R_row_index_65_scaled));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : array_obj_ref_62_index_0_scale array_obj_ref_67_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      data_in <= R_row_index_60_resized & R_row_index_65_resized;
      R_row_index_60_scaled <= data_out(13 downto 7);
      R_row_index_65_scaled <= data_out(6 downto 0);
      guard_vector(0)  <=  not read_write_bar_1_buffer(0);
      guard_vector(1)  <= read_write_bar_1_buffer(0);
      reqL_unguarded(1) <= array_obj_ref_62_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_67_index_0_scale_req_0;
      array_obj_ref_62_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_67_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= array_obj_ref_62_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_67_index_0_scale_req_1;
      array_obj_ref_62_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_67_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_0_accessRegulator_0: access_regulator_base generic map (name => "ApIntMul_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      ApIntMul_group_0_accessRegulator_1: access_regulator_base generic map (name => "ApIntMul_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      ApIntMul_group_0_gI: SplitGuardInterface generic map(name => "ApIntMul_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          name => "ApIntMul_group_0",
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0001000",
          constant_width => 7,
          use_constant  => true,
          full_rate  => false,
          no_arbitration => false,
          min_clock_period => false,
          num_reqs => 2,
          use_input_buffering => true,
          detailed_buffering_per_input => inBUFs,
          detailed_buffering_per_output => outBUFs --
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator array_obj_ref_62_index_sum_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_62_index_sum_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_sum_1:started:   inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_col_index_61_scaled = "& Convert_SLV_To_Hex_String(R_col_index_61_scaled) & " R_row_index_60_scaled = "& Convert_SLV_To_Hex_String(R_row_index_60_scaled));
          --
        end if; 
        if array_obj_ref_62_index_sum_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_index_sum_1:finished:  outputs: " & " array_obj_ref_62_index_partial_sum_1= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_index_partial_sum_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : array_obj_ref_62_index_sum_1 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_index_61_scaled & R_row_index_60_scaled;
      array_obj_ref_62_index_partial_sum_1 <= data_out(6 downto 0);
      guard_vector(0)  <= read_write_bar_1_buffer(0);
      reqL_unguarded(0) <= array_obj_ref_62_index_sum_1_req_0;
      array_obj_ref_62_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_62_index_sum_1_req_1;
      array_obj_ref_62_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 7, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator array_obj_ref_67_index_sum_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_67_index_sum_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_sum_1:started:   inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " R_col_index_66_scaled = "& Convert_SLV_To_Hex_String(R_col_index_66_scaled) & " R_row_index_65_scaled = "& Convert_SLV_To_Hex_String(R_row_index_65_scaled));
          --
        end if; 
        if array_obj_ref_67_index_sum_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_index_sum_1:finished:  outputs: " & " array_obj_ref_67_index_partial_sum_1= "  & Convert_SLV_To_Hex_String(array_obj_ref_67_index_partial_sum_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : array_obj_ref_67_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_index_66_scaled & R_row_index_65_scaled;
      array_obj_ref_67_index_partial_sum_1 <= data_out(6 downto 0);
      guard_vector(0)  <=  not read_write_bar_1_buffer(0);
      reqL_unguarded(0) <= array_obj_ref_67_index_sum_1_req_0;
      array_obj_ref_67_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_67_index_sum_1_req_1;
      array_obj_ref_67_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 7, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator array_obj_ref_62_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_62_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_load_0:started:   inputs: " & " read_write_bar_1_buffer (guard)= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_62_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_62_word_address_0));
          --
        end if; 
        if array_obj_ref_62_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_62_load_0:finished:  outputs: " & " array_obj_ref_62_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_62_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_62_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_62_load_0_req_0,
        array_obj_ref_62_load_0_ack_0,
        array_obj_ref_62_load_0_req_1,
        array_obj_ref_62_load_0_ack_1,
        "array_obj_ref_62_load_0",
        "memory_space_3" ,
        array_obj_ref_62_data_0,
        array_obj_ref_62_word_address_0,
        "array_obj_ref_62_data_0",
        "array_obj_ref_62_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_62_load_0_req_0;
      array_obj_ref_62_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_62_load_0_req_1;
      array_obj_ref_62_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_write_bar_1_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_62_word_address_0;
      array_obj_ref_62_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(15 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_67_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_67_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_store_0:started:   inputs: " & " read_write_bar_1_buffer (guard complement )= " & Convert_SLV_To_String(read_write_bar_1_buffer) & " array_obj_ref_67_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_67_word_address_0) & " array_obj_ref_67_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_67_data_0));
          --
        end if; 
        if array_obj_ref_67_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMem:DP:array_obj_ref_67_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_67_store_0_req_0,
      array_obj_ref_67_store_0_ack_0,
      array_obj_ref_67_store_0_req_1,
      array_obj_ref_67_store_0_ack_1,
      "array_obj_ref_67_store_0",
      "memory_space_3" ,
      array_obj_ref_67_data_0,
      array_obj_ref_67_word_address_0,
      "array_obj_ref_67_data_0",
      "array_obj_ref_67_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_67_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(6 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_67_store_0_req_0;
      array_obj_ref_67_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_67_store_0_req_1;
      array_obj_ref_67_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_write_bar_1_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_67_word_address_0;
      data_in <= array_obj_ref_67_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(15 downto 0),
          mtag => memory_space_3_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end accessMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity cal_col_to_be_replaced is -- 
  generic (tag_length : integer); 
  port ( -- 
    J : in  std_logic_vector(4 downto 0);
    col_to_be_replaced : in  std_logic_vector(1 downto 0);
    new_col_to_be_replaced : out  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity cal_col_to_be_replaced;
architecture cal_col_to_be_replaced_arch of cal_col_to_be_replaced is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 7)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 2)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal J_buffer :  std_logic_vector(4 downto 0);
  signal J_update_enable: Boolean;
  signal col_to_be_replaced_buffer :  std_logic_vector(1 downto 0);
  signal col_to_be_replaced_update_enable: Boolean;
  -- output port buffer signals
  signal new_col_to_be_replaced_buffer :  std_logic_vector(1 downto 0);
  signal new_col_to_be_replaced_update_enable: Boolean;
  signal cal_col_to_be_replaced_CP_2404_start: Boolean;
  signal cal_col_to_be_replaced_CP_2404_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal MUX_597_inst_req_0 : boolean;
  signal MUX_597_inst_ack_0 : boolean;
  signal MUX_597_inst_req_1 : boolean;
  signal MUX_597_inst_ack_1 : boolean;
  signal MUX_613_inst_req_0 : boolean;
  signal MUX_613_inst_ack_0 : boolean;
  signal MUX_613_inst_req_1 : boolean;
  signal MUX_613_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "cal_col_to_be_replaced_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 7) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(4 downto 0) <= J;
  J_buffer <= in_buffer_data_out(4 downto 0);
  in_buffer_data_in(6 downto 5) <= col_to_be_replaced;
  col_to_be_replaced_buffer <= in_buffer_data_out(6 downto 5);
  in_buffer_data_in(tag_length + 6 downto 7) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 6 downto 7);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  cal_col_to_be_replaced_CP_2404_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "cal_col_to_be_replaced_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 2) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(1 downto 0) <= new_col_to_be_replaced_buffer;
  new_col_to_be_replaced <= out_buffer_data_out(1 downto 0);
  out_buffer_data_in(tag_length + 1 downto 2) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 1 downto 2);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= cal_col_to_be_replaced_CP_2404_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= cal_col_to_be_replaced_CP_2404_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= cal_col_to_be_replaced_CP_2404_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,cal_col_to_be_replaced_CP_2404_start,"cal_col_to_be_replaced cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,cal_col_to_be_replaced_CP_2404_symbol, "cal_col_to_be_replaced cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  cal_col_to_be_replaced_CP_2404: Block -- control-path 
    signal cal_col_to_be_replaced_CP_2404_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    cal_col_to_be_replaced_CP_2404_elements(0) <= cal_col_to_be_replaced_CP_2404_start;
    cal_col_to_be_replaced_CP_2404_symbol <= cal_col_to_be_replaced_CP_2404_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/$entry
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_sample_start_
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_update_start_
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_start/$entry
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_start/req
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_complete/$entry
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_complete/req
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_update_start_
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_complete/$entry
      -- CP-element group 0: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_complete/req
      -- 
    -- logger for CP element group cal_col_to_be_replaced_CP_2404_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and cal_col_to_be_replaced_CP_2404_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:cal_col_to_be_replaced_CP_2404_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_597_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_597_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_613_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cal_col_to_be_replaced_CP_2404_elements(0), ack => MUX_597_inst_req_0); -- 
    req_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cal_col_to_be_replaced_CP_2404_elements(0), ack => MUX_597_inst_req_1); -- 
    req_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cal_col_to_be_replaced_CP_2404_elements(0), ack => MUX_613_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_sample_completed_
      -- CP-element group 1: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_start/$exit
      -- CP-element group 1: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_start/ack
      -- 
    -- logger for CP element group cal_col_to_be_replaced_CP_2404_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and cal_col_to_be_replaced_CP_2404_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:cal_col_to_be_replaced_CP_2404_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_597_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_597_inst_ack_0, ack => cal_col_to_be_replaced_CP_2404_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_update_completed_
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_complete/$exit
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_597_complete/ack
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_sample_start_
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_start/$entry
      -- CP-element group 2: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_start/req
      -- 
    -- logger for CP element group cal_col_to_be_replaced_CP_2404_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and cal_col_to_be_replaced_CP_2404_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:cal_col_to_be_replaced_CP_2404_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_597_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_613_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_597_inst_ack_1, ack => cal_col_to_be_replaced_CP_2404_elements(2)); -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => cal_col_to_be_replaced_CP_2404_elements(2), ack => MUX_613_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_sample_completed_
      -- CP-element group 3: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_start/$exit
      -- CP-element group 3: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_start/ack
      -- 
    -- logger for CP element group cal_col_to_be_replaced_CP_2404_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and cal_col_to_be_replaced_CP_2404_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:cal_col_to_be_replaced_CP_2404_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_613_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_613_inst_ack_0, ack => cal_col_to_be_replaced_CP_2404_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_586_to_assign_stmt_614/$exit
      -- CP-element group 4: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_update_completed_
      -- CP-element group 4: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_complete/$exit
      -- CP-element group 4: 	 assign_stmt_586_to_assign_stmt_614/MUX_613_complete/ack
      -- 
    -- logger for CP element group cal_col_to_be_replaced_CP_2404_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and cal_col_to_be_replaced_CP_2404_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:cal_col_to_be_replaced_CP_2404_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:cal_col_to_be_replaced:CP:MUX_613_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_613_inst_ack_1, ack => cal_col_to_be_replaced_CP_2404_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u2_u2_595_wire : std_logic_vector(1 downto 0);
    signal EQ_u2_u1_590_wire : std_logic_vector(0 downto 0);
    signal EQ_u5_u1_602_wire : std_logic_vector(0 downto 0);
    signal R_last_value_J_601_wire_constant : std_logic_vector(4 downto 0);
    signal checkJZero_608 : std_logic_vector(0 downto 0);
    signal col_to_be_replaced_3_586 : std_logic_vector(1 downto 0);
    signal col_to_be_replaced_other_598 : std_logic_vector(1 downto 0);
    signal konst_589_wire_constant : std_logic_vector(1 downto 0);
    signal konst_594_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_592_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_596_wire : std_logic_vector(1 downto 0);
    signal type_cast_604_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_last_value_J_601_wire_constant <= "00100";
    col_to_be_replaced_3_586 <= "11";
    konst_589_wire_constant <= "11";
    konst_594_wire_constant <= "01";
    type_cast_592_wire_constant <= "00";
    type_cast_604_wire_constant <= "0";
    type_cast_606_wire_constant <= "1";
    -- logger for split-operator MUX_597_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_597_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:MUX_597_inst:started:   inputs: " & " EQ_u2_u1_590_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_590_wire) & " type_cast_592_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_592_wire_constant) & " type_cast_596_wire = "& Convert_SLV_To_Hex_String(type_cast_596_wire));
          --
        end if; 
        if MUX_597_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:MUX_597_inst:finished:  outputs: " & " col_to_be_replaced_other_598= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_other_598));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_597_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_597_inst_req_0;
      MUX_597_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_597_inst_req_1;
      MUX_597_inst_ack_1<= update_ack(0);
      MUX_597_inst: SelectSplitProtocol generic map(name => "MUX_597_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_592_wire_constant, y => type_cast_596_wire, sel => EQ_u2_u1_590_wire, z => col_to_be_replaced_other_598, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_607_inst flow-through 
    process(checkJZero_608) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:MUX_607_inst:flowthrough inputs: " & " EQ_u5_u1_602_wire = "& Convert_SLV_To_Hex_String(EQ_u5_u1_602_wire) & " type_cast_604_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_604_wire_constant) & " type_cast_606_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_606_wire_constant) & " outputs:" & " checkJZero_608= "  & Convert_SLV_To_Hex_String(checkJZero_608));
      --
    end process; 
    -- flow-through select operator MUX_607_inst
    checkJZero_608 <= type_cast_604_wire_constant when (EQ_u5_u1_602_wire(0) /=  '0') else type_cast_606_wire_constant;
    -- logger for split-operator MUX_613_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_613_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:MUX_613_inst:started:   inputs: " & " checkJZero_608 = "& Convert_SLV_To_Hex_String(checkJZero_608) & " col_to_be_replaced_other_598 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_other_598) & " col_to_be_replaced_3_586 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_586));
          --
        end if; 
        if MUX_613_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:MUX_613_inst:finished:  outputs: " & " new_col_to_be_replaced_buffer= "  & Convert_SLV_To_Hex_String(new_col_to_be_replaced_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_613_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_613_inst_req_0;
      MUX_613_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_613_inst_req_1;
      MUX_613_inst_ack_1<= update_ack(0);
      MUX_613_inst: SelectSplitProtocol generic map(name => "MUX_613_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => col_to_be_replaced_other_598, y => col_to_be_replaced_3_586, sel => checkJZero_608, z => new_col_to_be_replaced_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator type_cast_596_inst flow-through 
    process(type_cast_596_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:type_cast_596_inst:flowthrough inputs: " & " ADD_u2_u2_595_wire = "& Convert_SLV_To_Hex_String(ADD_u2_u2_595_wire) & " outputs:" & " type_cast_596_wire= "  & Convert_SLV_To_Hex_String(type_cast_596_wire));
      --
    end process; 
    -- interlock type_cast_596_inst
    process(ADD_u2_u2_595_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := ADD_u2_u2_595_wire(1 downto 0);
      type_cast_596_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ADD_u2_u2_595_inst flow-through 
    process(ADD_u2_u2_595_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:ADD_u2_u2_595_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_594_wire_constant = "& Convert_SLV_To_Hex_String(konst_594_wire_constant) & " outputs:" & " ADD_u2_u2_595_wire= "  & Convert_SLV_To_Hex_String(ADD_u2_u2_595_wire));
      --
    end process; 
    -- binary operator ADD_u2_u2_595_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_to_be_replaced_buffer, konst_594_wire_constant, tmp_var);
      ADD_u2_u2_595_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_590_inst flow-through 
    process(EQ_u2_u1_590_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:EQ_u2_u1_590_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_589_wire_constant = "& Convert_SLV_To_Hex_String(konst_589_wire_constant) & " outputs:" & " EQ_u2_u1_590_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_590_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_590_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_to_be_replaced_buffer, konst_589_wire_constant, tmp_var);
      EQ_u2_u1_590_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u5_u1_602_inst flow-through 
    process(EQ_u5_u1_602_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:cal_col_to_be_replaced:DP:EQ_u5_u1_602_inst:flowthrough inputs: " & " J_buffer = "& Convert_SLV_To_Hex_String(J_buffer) & " R_last_value_J_601_wire_constant = "& Convert_SLV_To_Hex_String(R_last_value_J_601_wire_constant) & " outputs:" & " EQ_u5_u1_602_wire= "  & Convert_SLV_To_Hex_String(EQ_u5_u1_602_wire));
      --
    end process; 
    -- binary operator EQ_u5_u1_602_inst
    process(J_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_buffer, R_last_value_J_601_wire_constant, tmp_var);
      EQ_u5_u1_602_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end cal_col_to_be_replaced_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity initFilter is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_row_filter : in  std_logic_vector(5 downto 0);
    filter_initialized : out  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initFilter;
architecture initFilter_arch of initFilter is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 2)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_row_filter_buffer :  std_logic_vector(5 downto 0);
  signal start_row_filter_update_enable: Boolean;
  -- output port buffer signals
  signal filter_initialized_buffer :  std_logic_vector(1 downto 0);
  signal initFilter_CP_326_start: Boolean;
  signal initFilter_CP_326_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_J_174_delayed_7_0_175_inst_ack_0 : boolean;
  signal W_J_174_delayed_7_0_175_inst_ack_1 : boolean;
  signal W_J_174_delayed_7_0_175_inst_req_1 : boolean;
  signal array_obj_ref_180_store_0_ack_0 : boolean;
  signal array_obj_ref_180_store_0_req_0 : boolean;
  signal W_J_174_delayed_7_0_175_inst_req_0 : boolean;
  signal array_obj_ref_180_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_180_index_sum_1_req_1 : boolean;
  signal array_obj_ref_180_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_180_index_sum_1_req_0 : boolean;
  signal phi_stmt_123_req_1 : boolean;
  signal phi_stmt_123_req_0 : boolean;
  signal phi_stmt_123_ack_0 : boolean;
  signal array_obj_ref_180_store_0_ack_1 : boolean;
  signal array_obj_ref_180_store_0_req_1 : boolean;
  signal do_while_stmt_121_branch_ack_0 : boolean;
  signal array_obj_ref_180_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_180_index_0_scale_req_1 : boolean;
  signal array_obj_ref_180_index_0_scale_ack_0 : boolean;
  signal do_while_stmt_121_branch_ack_1 : boolean;
  signal array_obj_ref_180_index_0_scale_req_0 : boolean;
  signal do_while_stmt_121_branch_req_0 : boolean;
  signal n_ele_143_127_buf_req_0 : boolean;
  signal n_ele_143_127_buf_ack_0 : boolean;
  signal n_ele_143_127_buf_req_1 : boolean;
  signal n_ele_143_127_buf_ack_1 : boolean;
  signal phi_stmt_128_req_1 : boolean;
  signal phi_stmt_128_req_0 : boolean;
  signal phi_stmt_128_ack_0 : boolean;
  signal n_J_154_132_buf_req_0 : boolean;
  signal n_J_154_132_buf_ack_0 : boolean;
  signal n_J_154_132_buf_req_1 : boolean;
  signal n_J_154_132_buf_ack_1 : boolean;
  signal phi_stmt_133_req_1 : boolean;
  signal phi_stmt_133_req_0 : boolean;
  signal phi_stmt_133_ack_0 : boolean;
  signal n_I_165_137_buf_req_0 : boolean;
  signal n_I_165_137_buf_ack_0 : boolean;
  signal n_I_165_137_buf_req_1 : boolean;
  signal n_I_165_137_buf_ack_1 : boolean;
  signal call_stmt_171_call_req_0 : boolean;
  signal call_stmt_171_call_ack_0 : boolean;
  signal call_stmt_171_call_req_1 : boolean;
  signal call_stmt_171_call_ack_1 : boolean;
  signal W_I_173_delayed_7_0_172_inst_req_0 : boolean;
  signal W_I_173_delayed_7_0_172_inst_ack_0 : boolean;
  signal W_I_173_delayed_7_0_172_inst_req_1 : boolean;
  signal W_I_173_delayed_7_0_172_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initFilter_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= start_row_filter;
  start_row_filter_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initFilter_CP_326_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initFilter_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 2) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  filter_initialized_buffer <= "01";
  out_buffer_data_in(1 downto 0) <= filter_initialized_buffer;
  filter_initialized <= out_buffer_data_out(1 downto 0);
  out_buffer_data_in(tag_length + 1 downto 2) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 1 downto 2);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initFilter_CP_326_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initFilter_CP_326_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initFilter_CP_326_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,initFilter_CP_326_start,"initFilter cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,initFilter_CP_326_symbol, "initFilter cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initFilter_CP_326: Block -- control-path 
    signal initFilter_CP_326_elements: BooleanArray(99 downto 0);
    -- 
  begin -- 
    initFilter_CP_326_elements(0) <= initFilter_CP_326_start;
    initFilter_CP_326_symbol <= initFilter_CP_326_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_120/$entry
      -- CP-element group 0: 	 branch_block_stmt_120/branch_block_stmt_120__entry__
      -- CP-element group 0: 	 branch_block_stmt_120/do_while_stmt_121__entry__
      -- 
    -- logger for CP element group initFilter_CP_326_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	99 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_191/$exit
      -- CP-element group 1: 	 assign_stmt_191/$entry
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_120/$exit
      -- CP-element group 1: 	 branch_block_stmt_120/branch_block_stmt_120__exit__
      -- CP-element group 1: 	 branch_block_stmt_120/do_while_stmt_121__exit__
      -- 
    -- logger for CP element group initFilter_CP_326_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(1) <= initFilter_CP_326_elements(99);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_120/do_while_stmt_121/$entry
      -- CP-element group 2: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121__entry__
      -- 
    -- logger for CP element group initFilter_CP_326_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(2) <= initFilter_CP_326_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	99 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121__exit__
      -- 
    -- logger for CP element group initFilter_CP_326_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_120/do_while_stmt_121/loop_back
      -- 
    -- logger for CP element group initFilter_CP_326_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	97 
    -- CP-element group 5: 	98 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_120/do_while_stmt_121/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_120/do_while_stmt_121/condition_done
      -- CP-element group 5: 	 branch_block_stmt_120/do_while_stmt_121/loop_exit/$entry
      -- 
    -- logger for CP element group initFilter_CP_326_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(5) <= initFilter_CP_326_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	96 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_120/do_while_stmt_121/loop_body_done
      -- 
    -- logger for CP element group initFilter_CP_326_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(6) <= initFilter_CP_326_elements(96);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	38 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group initFilter_CP_326_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(7) <= initFilter_CP_326_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	40 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group initFilter_CP_326_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(8) <= initFilter_CP_326_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	86 
    -- CP-element group 9: 	90 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	95 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/loop_body_start
      -- 
    -- logger for CP element group initFilter_CP_326_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	95 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/condition_evaluated
      -- 
    -- logger for CP element group initFilter_CP_326_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:do_while_stmt_121_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(10), ack => do_while_stmt_121_branch_req_0); -- 
    initFilter_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(14) & initFilter_CP_326_elements(95);
      gj_initFilter_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	32 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	34 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_sample_start__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(15) & initFilter_CP_326_elements(51) & initFilter_CP_326_elements(32) & initFilter_CP_326_elements(14);
      gj_initFilter_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	32 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_sample_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(17) & initFilter_CP_326_elements(54) & initFilter_CP_326_elements(35);
      gj_initFilter_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	36 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(16) & initFilter_CP_326_elements(52) & initFilter_CP_326_elements(33);
      gj_initFilter_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	37 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(18) & initFilter_CP_326_elements(56) & initFilter_CP_326_elements(37);
      gj_initFilter_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_sample_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(12);
      gj_initFilter_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(18);
      gj_initFilter_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_sample_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_loopback_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(19) <= initFilter_CP_326_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_loopback_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_123_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_123_loopback_sample_req_365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_123_loopback_sample_req_365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(20), ack => phi_stmt_123_req_1); -- 
    -- Element group initFilter_CP_326_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_entry_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(21) <= initFilter_CP_326_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_entry_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_123_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_123_entry_sample_req_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_123_entry_sample_req_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(22), ack => phi_stmt_123_req_0); -- 
    -- Element group initFilter_CP_326_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_123_phi_mux_ack_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_123_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_123_phi_mux_ack_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_123_ack_0, ack => initFilter_CP_326_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_sample_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_update_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(26) <= initFilter_CP_326_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_126_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => initFilter_CP_326_elements(25), ack => initFilter_CP_326_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Sample/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_ele_143_127_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(28), ack => n_ele_143_127_buf_req_0); -- 
    -- Element group initFilter_CP_326_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_update_start_
      -- CP-element group 29: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Update/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_ele_143_127_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(29), ack => n_ele_143_127_buf_req_1); -- 
    -- Element group initFilter_CP_326_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Sample/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_ele_143_127_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_ele_143_127_buf_ack_0, ack => initFilter_CP_326_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_ele_127_Update/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_ele_143_127_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_ele_143_127_buf_ack_1, ack => initFilter_CP_326_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_sample_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(12);
      gj_initFilter_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	80 
    -- CP-element group 33: 	72 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(80) & initFilter_CP_326_elements(72);
      gj_initFilter_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_sample_start__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(34) <= initFilter_CP_326_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_sample_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_update_start__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(36) <= initFilter_CP_326_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	70 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_update_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_loopback_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(38) <= initFilter_CP_326_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_loopback_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_128_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_128_loopback_sample_req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_loopback_sample_req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(39), ack => phi_stmt_128_req_1); -- 
    -- Element group initFilter_CP_326_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_entry_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(40) <= initFilter_CP_326_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_entry_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_128_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_128_entry_sample_req_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_128_entry_sample_req_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(41), ack => phi_stmt_128_req_0); -- 
    -- Element group initFilter_CP_326_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_128_phi_mux_ack_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_128_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_128_phi_mux_ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_128_ack_0, ack => initFilter_CP_326_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_sample_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_update_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(45) <= initFilter_CP_326_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_131_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => initFilter_CP_326_elements(44), ack => initFilter_CP_326_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Sample/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_J_154_132_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(47), ack => n_J_154_132_buf_req_0); -- 
    -- Element group initFilter_CP_326_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_update_start_
      -- CP-element group 48: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Update/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_J_154_132_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(48), ack => n_J_154_132_buf_req_1); -- 
    -- Element group initFilter_CP_326_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Sample/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_J_154_132_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_J_154_132_buf_ack_0, ack => initFilter_CP_326_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_J_132_Update/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_J_154_132_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_J_154_132_buf_ack_1, ack => initFilter_CP_326_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_sample_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(12);
      gj_initFilter_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	76 
    -- CP-element group 52: 	72 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(52) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(76) & initFilter_CP_326_elements(72);
      gj_initFilter_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_sample_start__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(53) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(53) <= initFilter_CP_326_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_sample_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(54) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_update_start__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(55) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(55) <= initFilter_CP_326_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	74 
    -- CP-element group 56: 	70 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_update_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(56) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_loopback_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(57) <= initFilter_CP_326_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_loopback_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_133_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_133_loopback_sample_req_453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_loopback_sample_req_453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(58), ack => phi_stmt_133_req_1); -- 
    -- Element group initFilter_CP_326_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_entry_trigger
      -- 
    -- logger for CP element group initFilter_CP_326_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(59) <= initFilter_CP_326_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_entry_sample_req_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_133_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_133_entry_sample_req_456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_entry_sample_req_456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(60), ack => phi_stmt_133_req_0); -- 
    -- Element group initFilter_CP_326_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/phi_stmt_133_phi_mux_ack_ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:phi_stmt_133_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_133_phi_mux_ack_459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_133_ack_0, ack => initFilter_CP_326_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_sample_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(63) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_update_completed__ps
      -- 
    -- logger for CP element group initFilter_CP_326_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(64) <= initFilter_CP_326_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/type_cast_136_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => initFilter_CP_326_elements(63), ack => initFilter_CP_326_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Sample/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_I_165_137_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(66), ack => n_I_165_137_buf_req_0); -- 
    -- Element group initFilter_CP_326_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_update_start_
      -- CP-element group 67: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Update/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_I_165_137_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(67), ack => n_I_165_137_buf_req_1); -- 
    -- Element group initFilter_CP_326_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Sample/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_I_165_137_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_I_165_137_buf_ack_0, ack => initFilter_CP_326_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/R_n_I_137_Update/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:n_I_165_137_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_I_165_137_buf_ack_1, ack => initFilter_CP_326_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	56 
    -- CP-element group 70: 	37 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Sample/crr
      -- 
    -- logger for CP element group initFilter_CP_326_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:call_stmt_171_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(70), ack => call_stmt_171_call_req_0); -- 
    initFilter_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(56) & initFilter_CP_326_elements(37) & initFilter_CP_326_elements(72);
      gj_initFilter_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	93 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_update_start_
      -- CP-element group 71: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Update/ccr
      -- 
    -- logger for CP element group initFilter_CP_326_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:call_stmt_171_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(71), ack => call_stmt_171_call_req_1); -- 
    initFilter_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= initFilter_CP_326_elements(93);
      gj_initFilter_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	52 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	33 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Sample/cra
      -- 
    -- logger for CP element group initFilter_CP_326_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:call_stmt_171_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_171_call_ack_0, ack => initFilter_CP_326_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/call_stmt_171_Update/cca
      -- 
    -- logger for CP element group initFilter_CP_326_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:call_stmt_171_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_171_call_ack_1, ack => initFilter_CP_326_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	56 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Sample/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_I_173_delayed_7_0_172_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(74), ack => W_I_173_delayed_7_0_172_inst_req_0); -- 
    initFilter_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(56) & initFilter_CP_326_elements(76);
      gj_initFilter_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	84 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_update_start_
      -- CP-element group 75: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Update/req
      -- 
    -- logger for CP element group initFilter_CP_326_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_I_173_delayed_7_0_172_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(75), ack => W_I_173_delayed_7_0_172_inst_req_1); -- 
    initFilter_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(84) & initFilter_CP_326_elements(77);
      gj_initFilter_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	52 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Sample/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_I_173_delayed_7_0_172_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_173_delayed_7_0_172_inst_ack_0, ack => initFilter_CP_326_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_0/index_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_0/index_resize_req
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_computed_0
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resized_0
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_174_Update/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_I_173_delayed_7_0_172_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_I_173_delayed_7_0_172_inst_ack_1, ack => initFilter_CP_326_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Sample/req
      -- CP-element group 78: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_sample_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_J_174_delayed_7_0_175_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(78), ack => W_J_174_delayed_7_0_175_inst_req_0); -- 
    initFilter_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(37) & initFilter_CP_326_elements(80);
      gj_initFilter_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	91 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Update/req
      -- CP-element group 79: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_update_start_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_J_174_delayed_7_0_175_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(79), ack => W_J_174_delayed_7_0_175_inst_req_1); -- 
    initFilter_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= initFilter_CP_326_elements(91);
      gj_initFilter_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	33 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_sample_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_J_174_delayed_7_0_175_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_174_delayed_7_0_175_inst_ack_0, ack => initFilter_CP_326_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (14) 
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Update/ack
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_1/scale_rename_ack
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_1/scale_rename_req
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_1/$exit
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_1/$entry
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_1/index_resize_ack
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_1/index_resize_req
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_1/$exit
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resize_1/$entry
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_computed_1
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scaled_1
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_resized_1
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/assign_stmt_177_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:W_J_174_delayed_7_0_175_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_J_174_delayed_7_0_175_inst_ack_1, ack => initFilter_CP_326_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	92 
    -- CP-element group 82: 	73 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	93 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	93 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/word_0/rr
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/word_0/$entry
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/$entry
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/array_obj_ref_180_Split/split_ack
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/array_obj_ref_180_Split/split_req
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/array_obj_ref_180_Split/$exit
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/array_obj_ref_180_Split/$entry
      -- CP-element group 82: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/$entry
      -- 
    -- logger for CP element group initFilter_CP_326_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(82), ack => array_obj_ref_180_store_0_req_0); -- 
    initFilter_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(92) & initFilter_CP_326_elements(73) & initFilter_CP_326_elements(93);
      gj_initFilter_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	94 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	94 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_update_start_
      -- CP-element group 83: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/word_0/cr
      -- CP-element group 83: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/word_0/$entry
      -- CP-element group 83: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/$entry
      -- 
    -- logger for CP element group initFilter_CP_326_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(83), ack => array_obj_ref_180_store_0_req_1); -- 
    initFilter_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= initFilter_CP_326_elements(94);
      gj_initFilter_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	88 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	89 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	75 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scaled_0
      -- 
    -- logger for CP element group initFilter_CP_326_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(88) & initFilter_CP_326_elements(91);
      gj_initFilter_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	77 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_sample_start
      -- CP-element group 85: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Sample/$entry
      -- 
    -- logger for CP element group initFilter_CP_326_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_0_scale_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(85), ack => array_obj_ref_180_index_0_scale_req_0); -- 
    initFilter_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(77) & initFilter_CP_326_elements(87);
      gj_initFilter_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	9 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_update_start
      -- CP-element group 86: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Update/$entry
      -- 
    -- logger for CP element group initFilter_CP_326_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_0_scale_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(86), ack => array_obj_ref_180_index_0_scale_req_1); -- 
    initFilter_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(88);
      gj_initFilter_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	96 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Sample/$exit
      -- 
    -- logger for CP element group initFilter_CP_326_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_0_scale_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_index_0_scale_ack_0, ack => initFilter_CP_326_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_index_scale_0_update_complete
      -- 
    -- logger for CP element group initFilter_CP_326_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_0_scale_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_index_0_scale_ack_1, ack => initFilter_CP_326_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	84 
    -- CP-element group 89: 	81 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_sample_start
      -- 
    -- logger for CP element group initFilter_CP_326_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_sum_1_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(89), ack => array_obj_ref_180_index_sum_1_req_0); -- 
    initFilter_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(84) & initFilter_CP_326_elements(81) & initFilter_CP_326_elements(91);
      gj_initFilter_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	9 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	93 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_update_start
      -- 
    -- logger for CP element group initFilter_CP_326_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_sum_1_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initFilter_CP_326_elements(90), ack => array_obj_ref_180_index_sum_1_req_1); -- 
    initFilter_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(9) & initFilter_CP_326_elements(93);
      gj_initFilter_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	96 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	84 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	79 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_sample_complete
      -- 
    -- logger for CP element group initFilter_CP_326_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_sum_1_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_index_sum_1_ack_0, ack => initFilter_CP_326_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	82 
    -- CP-element group 92:  members (18) 
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_root_address_calculated
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_word_address_calculated
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_word_addrgen/root_register_ack
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_word_addrgen/root_register_req
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_word_addrgen/$exit
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_word_addrgen/$entry
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_base_plus_offset/sum_rename_ack
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_base_plus_offset/sum_rename_req
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_base_plus_offset/$exit
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_base_plus_offset/$entry
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_final_index_sum_regn/ack
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_final_index_sum_regn/req
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_final_index_sum_regn/$exit
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_final_index_sum_regn/$entry
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_partial_sum_1_update_complete
      -- CP-element group 92: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_offset_calculated
      -- 
    -- logger for CP element group initFilter_CP_326_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_index_sum_1_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_index_sum_1_ack_1, ack => initFilter_CP_326_elements(92)); -- 
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	82 
    -- CP-element group 93: successors 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: 	82 
    -- CP-element group 93: 	71 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/word_0/ra
      -- CP-element group 93: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/word_access_start/$exit
      -- CP-element group 93: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Sample/$exit
      -- 
    -- logger for CP element group initFilter_CP_326_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_store_0_ack_0, ack => initFilter_CP_326_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	83 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	83 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/word_access_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/array_obj_ref_180_update_completed_
      -- 
    -- logger for CP element group initFilter_CP_326_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:array_obj_ref_180_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_180_store_0_ack_1, ack => initFilter_CP_326_elements(94)); -- 
    -- CP-element group 95:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	9 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	10 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group initFilter_CP_326_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(95) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initFilter_CP_326_elements(95) is a control-delay.
    cp_element_95_delay: control_delay_element  generic map(name => " 95_delay", delay_value => 1)  port map(req => initFilter_CP_326_elements(9), ack => initFilter_CP_326_elements(95), clk => clk, reset =>reset);
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: 	87 
    -- CP-element group 96: 	91 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	6 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_120/do_while_stmt_121/do_while_stmt_121_loop_body/$exit
      -- 
    -- logger for CP element group initFilter_CP_326_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(96) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "initFilter_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= initFilter_CP_326_elements(12) & initFilter_CP_326_elements(87) & initFilter_CP_326_elements(91) & initFilter_CP_326_elements(94);
      gj_initFilter_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initFilter_CP_326_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	5 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_120/do_while_stmt_121/loop_exit/$exit
      -- CP-element group 97: 	 branch_block_stmt_120/do_while_stmt_121/loop_exit/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:do_while_stmt_121_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_121_branch_ack_0, ack => initFilter_CP_326_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	5 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_120/do_while_stmt_121/loop_taken/$exit
      -- CP-element group 98: 	 branch_block_stmt_120/do_while_stmt_121/loop_taken/ack
      -- 
    -- logger for CP element group initFilter_CP_326_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:do_while_stmt_121_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_121_branch_ack_1, ack => initFilter_CP_326_elements(98)); -- 
    -- CP-element group 99:  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	3 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	1 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_120/do_while_stmt_121/$exit
      -- 
    -- logger for CP element group initFilter_CP_326_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initFilter_CP_326_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initFilter:CP:initFilter_CP_326_elements(99) fired."); 
        -- 
      end if; --
    end process; 
    initFilter_CP_326_elements(99) <= initFilter_CP_326_elements(3);
    initFilter_do_while_stmt_121_terminator_637: loop_terminator -- 
      generic map (name => " initFilter_do_while_stmt_121_terminator_637", max_iterations_in_flight =>7) 
      port map(loop_body_exit => initFilter_CP_326_elements(6),loop_continue => initFilter_CP_326_elements(98),loop_terminate => initFilter_CP_326_elements(97),loop_back => initFilter_CP_326_elements(4),loop_exit => initFilter_CP_326_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_123_phi_seq_399_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initFilter_CP_326_elements(21);
      initFilter_CP_326_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initFilter_CP_326_elements(24);
      initFilter_CP_326_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= initFilter_CP_326_elements(26);
      initFilter_CP_326_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= initFilter_CP_326_elements(19);
      initFilter_CP_326_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initFilter_CP_326_elements(30);
      initFilter_CP_326_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= initFilter_CP_326_elements(31);
      initFilter_CP_326_elements(20) <= phi_mux_reqs(1);
      phi_stmt_123_phi_seq_399 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_123_phi_seq_399") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initFilter_CP_326_elements(11), 
          phi_sample_ack => initFilter_CP_326_elements(17), 
          phi_update_req => initFilter_CP_326_elements(13), 
          phi_update_ack => initFilter_CP_326_elements(18), 
          phi_mux_ack => initFilter_CP_326_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_128_phi_seq_443_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initFilter_CP_326_elements(40);
      initFilter_CP_326_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initFilter_CP_326_elements(43);
      initFilter_CP_326_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= initFilter_CP_326_elements(45);
      initFilter_CP_326_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= initFilter_CP_326_elements(38);
      initFilter_CP_326_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initFilter_CP_326_elements(49);
      initFilter_CP_326_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= initFilter_CP_326_elements(50);
      initFilter_CP_326_elements(39) <= phi_mux_reqs(1);
      phi_stmt_128_phi_seq_443 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_128_phi_seq_443") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initFilter_CP_326_elements(34), 
          phi_sample_ack => initFilter_CP_326_elements(35), 
          phi_update_req => initFilter_CP_326_elements(36), 
          phi_update_ack => initFilter_CP_326_elements(37), 
          phi_mux_ack => initFilter_CP_326_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_133_phi_seq_487_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= initFilter_CP_326_elements(59);
      initFilter_CP_326_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= initFilter_CP_326_elements(62);
      initFilter_CP_326_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= initFilter_CP_326_elements(64);
      initFilter_CP_326_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= initFilter_CP_326_elements(57);
      initFilter_CP_326_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= initFilter_CP_326_elements(68);
      initFilter_CP_326_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= initFilter_CP_326_elements(69);
      initFilter_CP_326_elements(58) <= phi_mux_reqs(1);
      phi_stmt_133_phi_seq_487 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_133_phi_seq_487") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => initFilter_CP_326_elements(53), 
          phi_sample_ack => initFilter_CP_326_elements(54), 
          phi_update_req => initFilter_CP_326_elements(55), 
          phi_update_ack => initFilter_CP_326_elements(56), 
          phi_mux_ack => initFilter_CP_326_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_351_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= initFilter_CP_326_elements(7);
        preds(1)  <= initFilter_CP_326_elements(8);
        entry_tmerge_351 : transition_merge -- 
          generic map(name => " entry_tmerge_351")
          port map (preds => preds, symbol_out => initFilter_CP_326_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_150_wire : std_logic_vector(4 downto 0);
    signal ADD_u6_u6_161_wire : std_logic_vector(5 downto 0);
    signal EQ_u5_u1_158_wire : std_logic_vector(0 downto 0);
    signal I_133 : std_logic_vector(5 downto 0);
    signal I_173_delayed_7_0_174 : std_logic_vector(5 downto 0);
    signal J_128 : std_logic_vector(4 downto 0);
    signal J_174_delayed_7_0_177 : std_logic_vector(4 downto 0);
    signal R_I_173_delayed_7_0_178_resized : std_logic_vector(3 downto 0);
    signal R_I_173_delayed_7_0_178_scaled : std_logic_vector(3 downto 0);
    signal R_J_174_delayed_7_0_179_resized : std_logic_vector(3 downto 0);
    signal R_J_174_delayed_7_0_179_scaled : std_logic_vector(3 downto 0);
    signal R_read_signal_166_wire_constant : std_logic_vector(0 downto 0);
    signal R_write_data_zero_169_wire_constant : std_logic_vector(15 downto 0);
    signal ULE_u5_u1_147_wire : std_logic_vector(0 downto 0);
    signal ULT_u5_u1_186_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_180_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_180_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_index_partial_sum_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_180_word_offset_0 : std_logic_vector(3 downto 0);
    signal ele_123 : std_logic_vector(4 downto 0);
    signal konst_141_wire_constant : std_logic_vector(4 downto 0);
    signal konst_146_wire_constant : std_logic_vector(4 downto 0);
    signal konst_149_wire_constant : std_logic_vector(4 downto 0);
    signal konst_157_wire_constant : std_logic_vector(4 downto 0);
    signal konst_160_wire_constant : std_logic_vector(5 downto 0);
    signal konst_185_wire_constant : std_logic_vector(4 downto 0);
    signal n_I_165 : std_logic_vector(5 downto 0);
    signal n_I_165_137_buffered : std_logic_vector(5 downto 0);
    signal n_J_154 : std_logic_vector(4 downto 0);
    signal n_J_154_132_buffered : std_logic_vector(4 downto 0);
    signal n_ele_143 : std_logic_vector(4 downto 0);
    signal n_ele_143_127_buffered : std_logic_vector(4 downto 0);
    signal rdata_171 : std_logic_vector(15 downto 0);
    signal type_cast_126_wire_constant : std_logic_vector(4 downto 0);
    signal type_cast_131_wire_constant : std_logic_vector(4 downto 0);
    signal type_cast_136_wire_constant : std_logic_vector(5 downto 0);
    signal type_cast_152_wire_constant : std_logic_vector(4 downto 0);
    signal type_cast_162_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    R_read_signal_166_wire_constant <= "1";
    R_write_data_zero_169_wire_constant <= "0000000000000000";
    array_obj_ref_180_offset_scale_factor_0 <= "0100";
    array_obj_ref_180_offset_scale_factor_1 <= "0001";
    array_obj_ref_180_resized_base_address <= "0000";
    array_obj_ref_180_word_offset_0 <= "0000";
    konst_141_wire_constant <= "00001";
    konst_146_wire_constant <= "00010";
    konst_149_wire_constant <= "00001";
    konst_157_wire_constant <= "00011";
    konst_160_wire_constant <= "000001";
    konst_185_wire_constant <= "01111";
    type_cast_126_wire_constant <= "00000";
    type_cast_131_wire_constant <= "00000";
    type_cast_136_wire_constant <= "001000";
    type_cast_152_wire_constant <= "00000";
    -- logger for phi phi_stmt_123
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_123_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_123:input-0 type_cast_126_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_126_wire_constant));
          --
        end if;
        if phi_stmt_123_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_123:input-1 n_ele_143_127_buffered= " & Convert_SLV_To_Hex_String(n_ele_143_127_buffered));
          --
        end if;
        if phi_stmt_123_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initFilter:DP:phi_stmt_123:sample-completed");
          --
        end if;
        if phi_stmt_123_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initFilter:DP:phi_stmt_123:output ele_123= " & Convert_SLV_To_Hex_String(ele_123));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_123: Block -- phi operator 
      signal idata: std_logic_vector(9 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_126_wire_constant & n_ele_143_127_buffered;
      req <= phi_stmt_123_req_0 & phi_stmt_123_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_123",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 5) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_123_ack_0,
          idata => idata,
          odata => ele_123,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_123
    -- logger for phi phi_stmt_128
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_128_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_128:input-0 type_cast_131_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_131_wire_constant));
          --
        end if;
        if phi_stmt_128_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_128:input-1 n_J_154_132_buffered= " & Convert_SLV_To_Hex_String(n_J_154_132_buffered));
          --
        end if;
        if phi_stmt_128_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initFilter:DP:phi_stmt_128:sample-completed");
          --
        end if;
        if phi_stmt_128_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initFilter:DP:phi_stmt_128:output J_128= " & Convert_SLV_To_Hex_String(J_128));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_128: Block -- phi operator 
      signal idata: std_logic_vector(9 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_131_wire_constant & n_J_154_132_buffered;
      req <= phi_stmt_128_req_0 & phi_stmt_128_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_128",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 5) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_128_ack_0,
          idata => idata,
          odata => J_128,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_128
    -- logger for phi phi_stmt_133
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_133_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_133:input-0 type_cast_136_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_136_wire_constant));
          --
        end if;
        if phi_stmt_133_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:initFilter:DP:phi_stmt_133:input-1 n_I_165_137_buffered= " & Convert_SLV_To_Hex_String(n_I_165_137_buffered));
          --
        end if;
        if phi_stmt_133_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:initFilter:DP:phi_stmt_133:sample-completed");
          --
        end if;
        if phi_stmt_133_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:initFilter:DP:phi_stmt_133:output I_133= " & Convert_SLV_To_Hex_String(I_133));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_133: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_136_wire_constant & n_I_165_137_buffered;
      req <= phi_stmt_133_req_0 & phi_stmt_133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_133",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_133_ack_0,
          idata => idata,
          odata => I_133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_133
    -- logger for split-operator MUX_153_inst flow-through 
    process(n_J_154) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:MUX_153_inst:flowthrough inputs: " & " ULE_u5_u1_147_wire = "& Convert_SLV_To_Hex_String(ULE_u5_u1_147_wire) & " ADD_u5_u5_150_wire = "& Convert_SLV_To_Hex_String(ADD_u5_u5_150_wire) & " type_cast_152_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_152_wire_constant) & " outputs:" & " n_J_154= "  & Convert_SLV_To_Hex_String(n_J_154));
      --
    end process; 
    -- flow-through select operator MUX_153_inst
    n_J_154 <= ADD_u5_u5_150_wire when (ULE_u5_u1_147_wire(0) /=  '0') else type_cast_152_wire_constant;
    -- logger for split-operator MUX_164_inst flow-through 
    process(n_I_165) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:MUX_164_inst:flowthrough inputs: " & " EQ_u5_u1_158_wire = "& Convert_SLV_To_Hex_String(EQ_u5_u1_158_wire) & " type_cast_162_wire = "& Convert_SLV_To_Hex_String(type_cast_162_wire) & " I_133 = "& Convert_SLV_To_Hex_String(I_133) & " outputs:" & " n_I_165= "  & Convert_SLV_To_Hex_String(n_I_165));
      --
    end process; 
    -- flow-through select operator MUX_164_inst
    n_I_165 <= type_cast_162_wire when (EQ_u5_u1_158_wire(0) /=  '0') else I_133;
    -- logger for split-operator W_I_173_delayed_7_0_172_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_I_173_delayed_7_0_172_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:W_I_173_delayed_7_0_172_inst:started:   inputs: " & " I_133 = "& Convert_SLV_To_Hex_String(I_133));
          --
        end if; 
        if W_I_173_delayed_7_0_172_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:W_I_173_delayed_7_0_172_inst:finished:  outputs: " & " I_173_delayed_7_0_174= "  & Convert_SLV_To_Hex_String(I_173_delayed_7_0_174));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_I_173_delayed_7_0_172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_I_173_delayed_7_0_172_inst_req_0;
      W_I_173_delayed_7_0_172_inst_ack_0<= wack(0);
      rreq(0) <= W_I_173_delayed_7_0_172_inst_req_1;
      W_I_173_delayed_7_0_172_inst_ack_1<= rack(0);
      W_I_173_delayed_7_0_172_inst : InterlockBuffer generic map ( -- 
        name => "W_I_173_delayed_7_0_172_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => I_173_delayed_7_0_174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator W_J_174_delayed_7_0_175_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_J_174_delayed_7_0_175_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:W_J_174_delayed_7_0_175_inst:started:   inputs: " & " J_128 = "& Convert_SLV_To_Hex_String(J_128));
          --
        end if; 
        if W_J_174_delayed_7_0_175_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:W_J_174_delayed_7_0_175_inst:finished:  outputs: " & " J_174_delayed_7_0_177= "  & Convert_SLV_To_Hex_String(J_174_delayed_7_0_177));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_J_174_delayed_7_0_175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_J_174_delayed_7_0_175_inst_req_0;
      W_J_174_delayed_7_0_175_inst_ack_0<= wack(0);
      rreq(0) <= W_J_174_delayed_7_0_175_inst_req_1;
      W_J_174_delayed_7_0_175_inst_ack_1<= rack(0);
      W_J_174_delayed_7_0_175_inst : InterlockBuffer generic map ( -- 
        name => "W_J_174_delayed_7_0_175_inst",
        buffer_size => 7,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => J_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => J_174_delayed_7_0_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_I_165_137_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_I_165_137_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_I_165_137_buf:started:   inputs: " & " n_I_165 = "& Convert_SLV_To_Hex_String(n_I_165));
          --
        end if; 
        if n_I_165_137_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_I_165_137_buf:finished:  outputs: " & " n_I_165_137_buffered= "  & Convert_SLV_To_Hex_String(n_I_165_137_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_I_165_137_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_I_165_137_buf_req_0;
      n_I_165_137_buf_ack_0<= wack(0);
      rreq(0) <= n_I_165_137_buf_req_1;
      n_I_165_137_buf_ack_1<= rack(0);
      n_I_165_137_buf : InterlockBuffer generic map ( -- 
        name => "n_I_165_137_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_I_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_I_165_137_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_J_154_132_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_J_154_132_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_J_154_132_buf:started:   inputs: " & " n_J_154 = "& Convert_SLV_To_Hex_String(n_J_154));
          --
        end if; 
        if n_J_154_132_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_J_154_132_buf:finished:  outputs: " & " n_J_154_132_buffered= "  & Convert_SLV_To_Hex_String(n_J_154_132_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_J_154_132_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_J_154_132_buf_req_0;
      n_J_154_132_buf_ack_0<= wack(0);
      rreq(0) <= n_J_154_132_buf_req_1;
      n_J_154_132_buf_ack_1<= rack(0);
      n_J_154_132_buf : InterlockBuffer generic map ( -- 
        name => "n_J_154_132_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_J_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_J_154_132_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_ele_143_127_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_ele_143_127_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_ele_143_127_buf:started:   inputs: " & " n_ele_143 = "& Convert_SLV_To_Hex_String(n_ele_143));
          --
        end if; 
        if n_ele_143_127_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:n_ele_143_127_buf:finished:  outputs: " & " n_ele_143_127_buffered= "  & Convert_SLV_To_Hex_String(n_ele_143_127_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_ele_143_127_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_ele_143_127_buf_req_0;
      n_ele_143_127_buf_ack_0<= wack(0);
      rreq(0) <= n_ele_143_127_buf_req_1;
      n_ele_143_127_buf_ack_1<= rack(0);
      n_ele_143_127_buf : InterlockBuffer generic map ( -- 
        name => "n_ele_143_127_buf",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  true ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_ele_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_ele_143_127_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_162_inst flow-through 
    process(type_cast_162_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:type_cast_162_inst:flowthrough inputs: " & " ADD_u6_u6_161_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_161_wire) & " outputs:" & " type_cast_162_wire= "  & Convert_SLV_To_Hex_String(type_cast_162_wire));
      --
    end process; 
    -- interlock type_cast_162_inst
    process(ADD_u6_u6_161_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_161_wire(5 downto 0);
      type_cast_162_wire <= tmp_var; -- 
    end process;
    -- logger for operator array_obj_ref_180_addr_0 flow-through 
    process(array_obj_ref_180_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_addr_0:flowthrough  inputs: " & " array_obj_ref_180_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_180_root_address) & "outputs: " & " array_obj_ref_180_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_180_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_180_addr_0
    process(array_obj_ref_180_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_180_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_180_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_gather_scatter flow-through 
    process(array_obj_ref_180_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_gather_scatter:flowthrough  inputs: " & " rdata_171 = "& Convert_SLV_To_Hex_String(rdata_171) & "outputs: " & " array_obj_ref_180_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_180_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_180_gather_scatter
    process(rdata_171) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_171;
      ov(15 downto 0) := iv;
      array_obj_ref_180_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_index_0_resize flow-through 
    process(R_I_173_delayed_7_0_178_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_0_resize:flowthrough  inputs: " & " I_173_delayed_7_0_174 = "& Convert_SLV_To_Hex_String(I_173_delayed_7_0_174) & "outputs: " & " R_I_173_delayed_7_0_178_resized= "  & Convert_SLV_To_Hex_String(R_I_173_delayed_7_0_178_resized));
      --
    end process; 
    -- equivalence array_obj_ref_180_index_0_resize
    process(I_173_delayed_7_0_174) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_173_delayed_7_0_174;
      ov := iv(3 downto 0);
      R_I_173_delayed_7_0_178_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_index_1_rename flow-through 
    process(R_J_174_delayed_7_0_179_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_1_rename:flowthrough  inputs: " & " R_J_174_delayed_7_0_179_resized = "& Convert_SLV_To_Hex_String(R_J_174_delayed_7_0_179_resized) & "outputs: " & " R_J_174_delayed_7_0_179_scaled= "  & Convert_SLV_To_Hex_String(R_J_174_delayed_7_0_179_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_180_index_1_rename
    process(R_J_174_delayed_7_0_179_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_J_174_delayed_7_0_179_resized;
      ov(3 downto 0) := iv;
      R_J_174_delayed_7_0_179_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_index_1_resize flow-through 
    process(R_J_174_delayed_7_0_179_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_1_resize:flowthrough  inputs: " & " J_174_delayed_7_0_177 = "& Convert_SLV_To_Hex_String(J_174_delayed_7_0_177) & "outputs: " & " R_J_174_delayed_7_0_179_resized= "  & Convert_SLV_To_Hex_String(R_J_174_delayed_7_0_179_resized));
      --
    end process; 
    -- equivalence array_obj_ref_180_index_1_resize
    process(J_174_delayed_7_0_177) --
      variable iv : std_logic_vector(4 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := J_174_delayed_7_0_177;
      ov := iv(3 downto 0);
      R_J_174_delayed_7_0_179_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_index_offset flow-through 
    process(array_obj_ref_180_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_offset:flowthrough  inputs: " & " array_obj_ref_180_index_partial_sum_1 = "& Convert_SLV_To_Hex_String(array_obj_ref_180_index_partial_sum_1) & "outputs: " & " array_obj_ref_180_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_180_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_180_index_offset
    process(array_obj_ref_180_index_partial_sum_1) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_180_index_partial_sum_1;
      ov(3 downto 0) := iv;
      array_obj_ref_180_final_offset <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_180_root_address_inst flow-through 
    process(array_obj_ref_180_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_root_address_inst:flowthrough  inputs: " & " array_obj_ref_180_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_180_final_offset) & "outputs: " & " array_obj_ref_180_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_180_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_180_root_address_inst
    process(array_obj_ref_180_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_180_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_180_root_address <= ov(3 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_121_branch_req_0," req0 do_while_stmt_121_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_121_branch_ack_0," ack0 do_while_stmt_121_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_121_branch_ack_1," ack1 do_while_stmt_121_branch");
    do_while_stmt_121_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u5_u1_186_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_121_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_121_branch_req_0,
          ack0 => do_while_stmt_121_branch_ack_0,
          ack1 => do_while_stmt_121_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u5_u5_142_inst flow-through 
    process(n_ele_143) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:ADD_u5_u5_142_inst:flowthrough inputs: " & " ele_123 = "& Convert_SLV_To_Hex_String(ele_123) & " konst_141_wire_constant = "& Convert_SLV_To_Hex_String(konst_141_wire_constant) & " outputs:" & " n_ele_143= "  & Convert_SLV_To_Hex_String(n_ele_143));
      --
    end process; 
    -- binary operator ADD_u5_u5_142_inst
    process(ele_123) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ele_123, konst_141_wire_constant, tmp_var);
      n_ele_143 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u5_u5_150_inst flow-through 
    process(ADD_u5_u5_150_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:ADD_u5_u5_150_inst:flowthrough inputs: " & " J_128 = "& Convert_SLV_To_Hex_String(J_128) & " konst_149_wire_constant = "& Convert_SLV_To_Hex_String(konst_149_wire_constant) & " outputs:" & " ADD_u5_u5_150_wire= "  & Convert_SLV_To_Hex_String(ADD_u5_u5_150_wire));
      --
    end process; 
    -- binary operator ADD_u5_u5_150_inst
    process(J_128) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntAdd_proc(J_128, konst_149_wire_constant, tmp_var);
      ADD_u5_u5_150_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_161_inst flow-through 
    process(ADD_u6_u6_161_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:ADD_u6_u6_161_inst:flowthrough inputs: " & " I_133 = "& Convert_SLV_To_Hex_String(I_133) & " konst_160_wire_constant = "& Convert_SLV_To_Hex_String(konst_160_wire_constant) & " outputs:" & " ADD_u6_u6_161_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_161_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_161_inst
    process(I_133) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_133, konst_160_wire_constant, tmp_var);
      ADD_u6_u6_161_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u5_u1_158_inst flow-through 
    process(EQ_u5_u1_158_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:EQ_u5_u1_158_inst:flowthrough inputs: " & " J_128 = "& Convert_SLV_To_Hex_String(J_128) & " konst_157_wire_constant = "& Convert_SLV_To_Hex_String(konst_157_wire_constant) & " outputs:" & " EQ_u5_u1_158_wire= "  & Convert_SLV_To_Hex_String(EQ_u5_u1_158_wire));
      --
    end process; 
    -- binary operator EQ_u5_u1_158_inst
    process(J_128) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_128, konst_157_wire_constant, tmp_var);
      EQ_u5_u1_158_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULE_u5_u1_147_inst flow-through 
    process(ULE_u5_u1_147_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:ULE_u5_u1_147_inst:flowthrough inputs: " & " J_128 = "& Convert_SLV_To_Hex_String(J_128) & " konst_146_wire_constant = "& Convert_SLV_To_Hex_String(konst_146_wire_constant) & " outputs:" & " ULE_u5_u1_147_wire= "  & Convert_SLV_To_Hex_String(ULE_u5_u1_147_wire));
      --
    end process; 
    -- binary operator ULE_u5_u1_147_inst
    process(J_128) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(J_128, konst_146_wire_constant, tmp_var);
      ULE_u5_u1_147_wire <= tmp_var; --
    end process;
    -- logger for split-operator ULT_u5_u1_186_inst flow-through 
    process(ULT_u5_u1_186_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:ULT_u5_u1_186_inst:flowthrough inputs: " & " ele_123 = "& Convert_SLV_To_Hex_String(ele_123) & " konst_185_wire_constant = "& Convert_SLV_To_Hex_String(konst_185_wire_constant) & " outputs:" & " ULT_u5_u1_186_wire= "  & Convert_SLV_To_Hex_String(ULT_u5_u1_186_wire));
      --
    end process; 
    -- binary operator ULT_u5_u1_186_inst
    process(ele_123) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(ele_123, konst_185_wire_constant, tmp_var);
      ULT_u5_u1_186_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_180_index_0_scale
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_180_index_0_scale_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_0_scale:started:   inputs: " & " R_I_173_delayed_7_0_178_resized = "& Convert_SLV_To_Hex_String(R_I_173_delayed_7_0_178_resized) & " array_obj_ref_180_offset_scale_factor_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_180_offset_scale_factor_0));
          --
        end if; 
        if array_obj_ref_180_index_0_scale_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_0_scale:finished:  outputs: " & " R_I_173_delayed_7_0_178_scaled= "  & Convert_SLV_To_Hex_String(R_I_173_delayed_7_0_178_scaled));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (6) : array_obj_ref_180_index_0_scale 
    ApIntMul_group_6: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_I_173_delayed_7_0_178_resized;
      R_I_173_delayed_7_0_178_scaled <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_180_index_0_scale_req_0;
      array_obj_ref_180_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_180_index_0_scale_req_1;
      array_obj_ref_180_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_6_gI: SplitGuardInterface generic map(name => "ApIntMul_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- logger for split-operator array_obj_ref_180_index_sum_1
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_180_index_sum_1_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_sum_1:started:   inputs: " & " R_J_174_delayed_7_0_179_scaled = "& Convert_SLV_To_Hex_String(R_J_174_delayed_7_0_179_scaled) & " R_I_173_delayed_7_0_178_scaled = "& Convert_SLV_To_Hex_String(R_I_173_delayed_7_0_178_scaled));
          --
        end if; 
        if array_obj_ref_180_index_sum_1_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_index_sum_1:finished:  outputs: " & " array_obj_ref_180_index_partial_sum_1= "  & Convert_SLV_To_Hex_String(array_obj_ref_180_index_partial_sum_1));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (7) : array_obj_ref_180_index_sum_1 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_J_174_delayed_7_0_179_scaled & R_I_173_delayed_7_0_178_scaled;
      array_obj_ref_180_index_partial_sum_1 <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_180_index_sum_1_req_0;
      array_obj_ref_180_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_180_index_sum_1_req_1;
      array_obj_ref_180_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 4, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- logger for split-operator array_obj_ref_180_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_180_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_store_0:started:   inputs: " & " array_obj_ref_180_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_180_word_address_0) & " array_obj_ref_180_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_180_data_0));
          --
        end if; 
        if array_obj_ref_180_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:array_obj_ref_180_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_180_store_0_req_0,
      array_obj_ref_180_store_0_ack_0,
      array_obj_ref_180_store_0_req_1,
      array_obj_ref_180_store_0_ack_1,
      "array_obj_ref_180_store_0",
      "memory_space_0" ,
      array_obj_ref_180_data_0,
      array_obj_ref_180_word_address_0,
      "array_obj_ref_180_data_0",
      "array_obj_ref_180_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_180_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 7);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_180_store_0_req_0;
      array_obj_ref_180_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_180_store_0_req_1;
      array_obj_ref_180_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_180_word_address_0;
      data_in <= array_obj_ref_180_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(3 downto 0),
          mdata => memory_space_0_sr_data(15 downto 0),
          mtag => memory_space_0_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator call_stmt_171_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_171_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:call_stmt_171_call:started:  Call to module accessMem inputs: " & " R_read_signal_166_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_166_wire_constant) & " I_133 = "& Convert_SLV_To_Hex_String(I_133) & " J_128 = "& Convert_SLV_To_Hex_String(J_128) & " R_write_data_zero_169_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_169_wire_constant));
          --
        end if; 
        if call_stmt_171_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initFilter:DP:call_stmt_171_call:finished:  outputs: " & " rdata_171= "  & Convert_SLV_To_Hex_String(rdata_171));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_171_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_171_call_req_0;
      call_stmt_171_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_171_call_req_1;
      call_stmt_171_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_read_signal_166_wire_constant & I_133 & J_128 & R_write_data_zero_169_wire_constant;
      rdata_171 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 28,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 5,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end initFilter_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity initIfMaps is -- 
  generic (tag_length : integer); 
  port ( -- 
    start : in  std_logic_vector(0 downto 0);
    I : in  std_logic_vector(5 downto 0);
    J : in  std_logic_vector(4 downto 0);
    col_to_be_replaced : in  std_logic_vector(1 downto 0);
    finished : out  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity initIfMaps;
architecture initIfMaps_arch of initIfMaps is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 14)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 2)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_buffer :  std_logic_vector(0 downto 0);
  signal start_update_enable: Boolean;
  signal I_buffer :  std_logic_vector(5 downto 0);
  signal I_update_enable: Boolean;
  signal J_buffer :  std_logic_vector(4 downto 0);
  signal J_update_enable: Boolean;
  signal col_to_be_replaced_buffer :  std_logic_vector(1 downto 0);
  signal col_to_be_replaced_update_enable: Boolean;
  -- output port buffer signals
  signal finished_buffer :  std_logic_vector(1 downto 0);
  signal initIfMaps_CP_641_start: Boolean;
  signal initIfMaps_CP_641_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal array_obj_ref_393_store_0_req_0 : boolean;
  signal type_cast_223_inst_req_1 : boolean;
  signal type_cast_223_inst_ack_1 : boolean;
  signal array_obj_ref_482_store_0_ack_0 : boolean;
  signal array_obj_ref_399_store_0_ack_1 : boolean;
  signal array_obj_ref_399_store_0_req_1 : boolean;
  signal type_cast_211_inst_ack_1 : boolean;
  signal array_obj_ref_469_store_0_req_1 : boolean;
  signal type_cast_211_inst_req_1 : boolean;
  signal type_cast_229_inst_req_1 : boolean;
  signal type_cast_229_inst_req_0 : boolean;
  signal type_cast_229_inst_ack_0 : boolean;
  signal type_cast_229_inst_ack_1 : boolean;
  signal array_obj_ref_482_store_0_req_0 : boolean;
  signal call_stmt_465_call_req_0 : boolean;
  signal call_stmt_465_call_ack_1 : boolean;
  signal call_stmt_446_call_ack_1 : boolean;
  signal call_stmt_408_call_req_1 : boolean;
  signal array_obj_ref_399_store_0_req_0 : boolean;
  signal call_stmt_478_call_req_0 : boolean;
  signal array_obj_ref_469_store_0_req_0 : boolean;
  signal array_obj_ref_456_store_0_req_1 : boolean;
  signal call_stmt_465_call_ack_0 : boolean;
  signal call_stmt_491_call_req_1 : boolean;
  signal call_stmt_491_call_ack_1 : boolean;
  signal array_obj_ref_437_store_0_ack_0 : boolean;
  signal call_stmt_446_call_req_0 : boolean;
  signal array_obj_ref_450_store_0_req_0 : boolean;
  signal array_obj_ref_393_store_0_req_1 : boolean;
  signal array_obj_ref_469_store_0_ack_0 : boolean;
  signal call_stmt_465_call_req_1 : boolean;
  signal call_stmt_446_call_ack_0 : boolean;
  signal type_cast_223_inst_req_0 : boolean;
  signal type_cast_223_inst_ack_0 : boolean;
  signal array_obj_ref_393_store_0_ack_1 : boolean;
  signal call_stmt_478_call_ack_1 : boolean;
  signal call_stmt_408_call_req_0 : boolean;
  signal call_stmt_478_call_ack_0 : boolean;
  signal array_obj_ref_393_store_0_ack_0 : boolean;
  signal type_cast_211_inst_ack_0 : boolean;
  signal type_cast_211_inst_req_0 : boolean;
  signal type_cast_217_inst_ack_0 : boolean;
  signal call_stmt_491_call_req_0 : boolean;
  signal call_stmt_491_call_ack_0 : boolean;
  signal array_obj_ref_437_store_0_req_0 : boolean;
  signal type_cast_217_inst_ack_1 : boolean;
  signal call_stmt_446_call_req_1 : boolean;
  signal array_obj_ref_482_store_0_ack_1 : boolean;
  signal call_stmt_427_call_ack_1 : boolean;
  signal call_stmt_427_call_req_1 : boolean;
  signal call_stmt_268_call_req_0 : boolean;
  signal call_stmt_268_call_ack_0 : boolean;
  signal call_stmt_268_call_req_1 : boolean;
  signal call_stmt_268_call_ack_1 : boolean;
  signal call_stmt_255_call_ack_1 : boolean;
  signal array_obj_ref_450_store_0_req_1 : boolean;
  signal array_obj_ref_259_store_0_req_0 : boolean;
  signal array_obj_ref_259_store_0_ack_0 : boolean;
  signal call_stmt_427_call_ack_0 : boolean;
  signal call_stmt_427_call_req_0 : boolean;
  signal array_obj_ref_259_store_0_req_1 : boolean;
  signal array_obj_ref_259_store_0_ack_1 : boolean;
  signal array_obj_ref_495_store_0_ack_0 : boolean;
  signal array_obj_ref_456_store_0_ack_0 : boolean;
  signal type_cast_235_inst_ack_1 : boolean;
  signal array_obj_ref_437_store_0_req_1 : boolean;
  signal type_cast_235_inst_req_1 : boolean;
  signal array_obj_ref_431_store_0_ack_1 : boolean;
  signal array_obj_ref_456_store_0_ack_1 : boolean;
  signal type_cast_217_inst_req_0 : boolean;
  signal array_obj_ref_399_store_0_ack_0 : boolean;
  signal array_obj_ref_469_store_0_ack_1 : boolean;
  signal type_cast_217_inst_req_1 : boolean;
  signal array_obj_ref_482_store_0_req_1 : boolean;
  signal call_stmt_255_call_req_0 : boolean;
  signal call_stmt_255_call_ack_0 : boolean;
  signal call_stmt_255_call_req_1 : boolean;
  signal array_obj_ref_450_store_0_ack_1 : boolean;
  signal type_cast_235_inst_req_0 : boolean;
  signal type_cast_235_inst_ack_0 : boolean;
  signal array_obj_ref_437_store_0_ack_1 : boolean;
  signal call_stmt_478_call_req_1 : boolean;
  signal call_stmt_408_call_ack_0 : boolean;
  signal array_obj_ref_450_store_0_ack_0 : boolean;
  signal array_obj_ref_418_store_0_ack_1 : boolean;
  signal array_obj_ref_272_store_0_req_0 : boolean;
  signal array_obj_ref_272_store_0_ack_0 : boolean;
  signal array_obj_ref_418_store_0_req_1 : boolean;
  signal array_obj_ref_272_store_0_req_1 : boolean;
  signal array_obj_ref_272_store_0_ack_1 : boolean;
  signal array_obj_ref_456_store_0_req_0 : boolean;
  signal call_stmt_281_call_req_0 : boolean;
  signal call_stmt_281_call_ack_0 : boolean;
  signal call_stmt_281_call_req_1 : boolean;
  signal call_stmt_281_call_ack_1 : boolean;
  signal array_obj_ref_495_store_0_req_0 : boolean;
  signal array_obj_ref_418_store_0_ack_0 : boolean;
  signal array_obj_ref_418_store_0_req_0 : boolean;
  signal array_obj_ref_285_store_0_req_0 : boolean;
  signal array_obj_ref_285_store_0_ack_0 : boolean;
  signal array_obj_ref_285_store_0_req_1 : boolean;
  signal array_obj_ref_285_store_0_ack_1 : boolean;
  signal array_obj_ref_431_store_0_req_1 : boolean;
  signal call_stmt_294_call_req_0 : boolean;
  signal call_stmt_294_call_ack_0 : boolean;
  signal call_stmt_294_call_req_1 : boolean;
  signal call_stmt_294_call_ack_1 : boolean;
  signal array_obj_ref_298_store_0_req_0 : boolean;
  signal array_obj_ref_298_store_0_ack_0 : boolean;
  signal array_obj_ref_298_store_0_req_1 : boolean;
  signal array_obj_ref_298_store_0_ack_1 : boolean;
  signal array_obj_ref_304_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_ack_0 : boolean;
  signal array_obj_ref_412_store_0_ack_1 : boolean;
  signal array_obj_ref_412_store_0_req_1 : boolean;
  signal array_obj_ref_304_store_0_req_1 : boolean;
  signal array_obj_ref_304_store_0_ack_1 : boolean;
  signal call_stmt_313_call_req_0 : boolean;
  signal call_stmt_313_call_ack_0 : boolean;
  signal call_stmt_313_call_req_1 : boolean;
  signal call_stmt_313_call_ack_1 : boolean;
  signal array_obj_ref_412_store_0_ack_0 : boolean;
  signal array_obj_ref_317_store_0_req_0 : boolean;
  signal array_obj_ref_317_store_0_ack_0 : boolean;
  signal array_obj_ref_412_store_0_req_0 : boolean;
  signal array_obj_ref_317_store_0_req_1 : boolean;
  signal array_obj_ref_317_store_0_ack_1 : boolean;
  signal array_obj_ref_431_store_0_ack_0 : boolean;
  signal array_obj_ref_323_store_0_req_0 : boolean;
  signal array_obj_ref_323_store_0_ack_0 : boolean;
  signal array_obj_ref_323_store_0_req_1 : boolean;
  signal array_obj_ref_323_store_0_ack_1 : boolean;
  signal array_obj_ref_431_store_0_req_0 : boolean;
  signal call_stmt_332_call_req_0 : boolean;
  signal call_stmt_332_call_ack_0 : boolean;
  signal call_stmt_332_call_req_1 : boolean;
  signal call_stmt_332_call_ack_1 : boolean;
  signal array_obj_ref_336_store_0_req_0 : boolean;
  signal array_obj_ref_336_store_0_ack_0 : boolean;
  signal call_stmt_408_call_ack_1 : boolean;
  signal array_obj_ref_336_store_0_req_1 : boolean;
  signal array_obj_ref_336_store_0_ack_1 : boolean;
  signal array_obj_ref_342_store_0_req_0 : boolean;
  signal array_obj_ref_342_store_0_ack_0 : boolean;
  signal array_obj_ref_342_store_0_req_1 : boolean;
  signal array_obj_ref_342_store_0_ack_1 : boolean;
  signal call_stmt_351_call_req_0 : boolean;
  signal call_stmt_351_call_ack_0 : boolean;
  signal call_stmt_351_call_req_1 : boolean;
  signal call_stmt_351_call_ack_1 : boolean;
  signal array_obj_ref_355_store_0_req_0 : boolean;
  signal array_obj_ref_355_store_0_ack_0 : boolean;
  signal array_obj_ref_355_store_0_req_1 : boolean;
  signal array_obj_ref_355_store_0_ack_1 : boolean;
  signal array_obj_ref_361_store_0_req_0 : boolean;
  signal array_obj_ref_361_store_0_ack_0 : boolean;
  signal array_obj_ref_361_store_0_req_1 : boolean;
  signal array_obj_ref_361_store_0_ack_1 : boolean;
  signal call_stmt_370_call_req_0 : boolean;
  signal call_stmt_370_call_ack_0 : boolean;
  signal call_stmt_370_call_req_1 : boolean;
  signal call_stmt_370_call_ack_1 : boolean;
  signal array_obj_ref_374_store_0_req_0 : boolean;
  signal array_obj_ref_374_store_0_ack_0 : boolean;
  signal array_obj_ref_374_store_0_req_1 : boolean;
  signal array_obj_ref_374_store_0_ack_1 : boolean;
  signal array_obj_ref_380_store_0_req_0 : boolean;
  signal array_obj_ref_380_store_0_ack_0 : boolean;
  signal array_obj_ref_380_store_0_req_1 : boolean;
  signal array_obj_ref_380_store_0_ack_1 : boolean;
  signal call_stmt_389_call_req_0 : boolean;
  signal call_stmt_389_call_ack_0 : boolean;
  signal call_stmt_389_call_req_1 : boolean;
  signal call_stmt_389_call_ack_1 : boolean;
  signal array_obj_ref_495_store_0_req_1 : boolean;
  signal array_obj_ref_495_store_0_ack_1 : boolean;
  signal type_cast_502_inst_req_0 : boolean;
  signal type_cast_502_inst_ack_0 : boolean;
  signal type_cast_502_inst_req_1 : boolean;
  signal type_cast_502_inst_ack_1 : boolean;
  signal call_stmt_509_call_req_0 : boolean;
  signal call_stmt_509_call_ack_0 : boolean;
  signal call_stmt_509_call_req_1 : boolean;
  signal call_stmt_509_call_ack_1 : boolean;
  signal array_obj_ref_512_index_offset_req_0 : boolean;
  signal array_obj_ref_512_index_offset_ack_0 : boolean;
  signal array_obj_ref_512_index_offset_req_1 : boolean;
  signal array_obj_ref_512_index_offset_ack_1 : boolean;
  signal array_obj_ref_512_store_0_req_0 : boolean;
  signal array_obj_ref_512_store_0_ack_0 : boolean;
  signal array_obj_ref_512_store_0_req_1 : boolean;
  signal array_obj_ref_512_store_0_ack_1 : boolean;
  signal call_stmt_520_call_req_0 : boolean;
  signal call_stmt_520_call_ack_0 : boolean;
  signal call_stmt_520_call_req_1 : boolean;
  signal call_stmt_520_call_ack_1 : boolean;
  signal array_obj_ref_523_index_offset_req_0 : boolean;
  signal array_obj_ref_523_index_offset_ack_0 : boolean;
  signal array_obj_ref_523_index_offset_req_1 : boolean;
  signal array_obj_ref_523_index_offset_ack_1 : boolean;
  signal array_obj_ref_523_store_0_req_0 : boolean;
  signal array_obj_ref_523_store_0_ack_0 : boolean;
  signal array_obj_ref_523_store_0_req_1 : boolean;
  signal array_obj_ref_523_store_0_ack_1 : boolean;
  signal array_obj_ref_528_index_offset_req_0 : boolean;
  signal array_obj_ref_528_index_offset_ack_0 : boolean;
  signal array_obj_ref_528_index_offset_req_1 : boolean;
  signal array_obj_ref_528_index_offset_ack_1 : boolean;
  signal array_obj_ref_528_store_0_req_0 : boolean;
  signal array_obj_ref_528_store_0_ack_0 : boolean;
  signal array_obj_ref_528_store_0_req_1 : boolean;
  signal array_obj_ref_528_store_0_ack_1 : boolean;
  signal call_stmt_536_call_req_0 : boolean;
  signal call_stmt_536_call_ack_0 : boolean;
  signal call_stmt_536_call_req_1 : boolean;
  signal call_stmt_536_call_ack_1 : boolean;
  signal array_obj_ref_539_index_offset_req_0 : boolean;
  signal array_obj_ref_539_index_offset_ack_0 : boolean;
  signal array_obj_ref_539_index_offset_req_1 : boolean;
  signal array_obj_ref_539_index_offset_ack_1 : boolean;
  signal array_obj_ref_539_store_0_req_0 : boolean;
  signal array_obj_ref_539_store_0_ack_0 : boolean;
  signal array_obj_ref_539_store_0_req_1 : boolean;
  signal array_obj_ref_539_store_0_ack_1 : boolean;
  signal array_obj_ref_544_index_offset_req_0 : boolean;
  signal array_obj_ref_544_index_offset_ack_0 : boolean;
  signal array_obj_ref_544_index_offset_req_1 : boolean;
  signal array_obj_ref_544_index_offset_ack_1 : boolean;
  signal array_obj_ref_544_store_0_req_0 : boolean;
  signal array_obj_ref_544_store_0_ack_0 : boolean;
  signal array_obj_ref_544_store_0_req_1 : boolean;
  signal array_obj_ref_544_store_0_ack_1 : boolean;
  signal call_stmt_552_call_req_0 : boolean;
  signal call_stmt_552_call_ack_0 : boolean;
  signal call_stmt_552_call_req_1 : boolean;
  signal call_stmt_552_call_ack_1 : boolean;
  signal array_obj_ref_555_index_offset_req_0 : boolean;
  signal array_obj_ref_555_index_offset_ack_0 : boolean;
  signal array_obj_ref_555_index_offset_req_1 : boolean;
  signal array_obj_ref_555_index_offset_ack_1 : boolean;
  signal array_obj_ref_555_store_0_req_0 : boolean;
  signal array_obj_ref_555_store_0_ack_0 : boolean;
  signal array_obj_ref_555_store_0_req_1 : boolean;
  signal array_obj_ref_555_store_0_ack_1 : boolean;
  signal array_obj_ref_560_index_offset_req_0 : boolean;
  signal array_obj_ref_560_index_offset_ack_0 : boolean;
  signal array_obj_ref_560_index_offset_req_1 : boolean;
  signal array_obj_ref_560_index_offset_ack_1 : boolean;
  signal array_obj_ref_560_store_0_req_0 : boolean;
  signal array_obj_ref_560_store_0_ack_0 : boolean;
  signal array_obj_ref_560_store_0_req_1 : boolean;
  signal array_obj_ref_560_store_0_ack_1 : boolean;
  signal call_stmt_568_call_req_0 : boolean;
  signal call_stmt_568_call_ack_0 : boolean;
  signal call_stmt_568_call_req_1 : boolean;
  signal call_stmt_568_call_ack_1 : boolean;
  signal array_obj_ref_571_index_offset_req_0 : boolean;
  signal array_obj_ref_571_index_offset_ack_0 : boolean;
  signal array_obj_ref_571_index_offset_req_1 : boolean;
  signal array_obj_ref_571_index_offset_ack_1 : boolean;
  signal array_obj_ref_571_store_0_req_0 : boolean;
  signal array_obj_ref_571_store_0_ack_0 : boolean;
  signal array_obj_ref_571_store_0_req_1 : boolean;
  signal array_obj_ref_571_store_0_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "initIfMaps_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 14) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= start;
  start_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(6 downto 1) <= I;
  I_buffer <= in_buffer_data_out(6 downto 1);
  in_buffer_data_in(11 downto 7) <= J;
  J_buffer <= in_buffer_data_out(11 downto 7);
  in_buffer_data_in(13 downto 12) <= col_to_be_replaced;
  col_to_be_replaced_buffer <= in_buffer_data_out(13 downto 12);
  in_buffer_data_in(tag_length + 13 downto 14) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 13 downto 14);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  initIfMaps_CP_641_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "initIfMaps_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 2) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  finished_buffer <= "01";
  out_buffer_data_in(1 downto 0) <= finished_buffer;
  finished <= out_buffer_data_out(1 downto 0);
  out_buffer_data_in(tag_length + 1 downto 2) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 1 downto 2);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initIfMaps_CP_641_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= initIfMaps_CP_641_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= initIfMaps_CP_641_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,initIfMaps_CP_641_start,"initIfMaps cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,initIfMaps_CP_641_symbol, "initIfMaps cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  initIfMaps_CP_641: Block -- control-path 
    signal initIfMaps_CP_641_elements: BooleanArray(233 downto 0);
    -- 
  begin -- 
    initIfMaps_CP_641_elements(0) <= initIfMaps_CP_641_start;
    initIfMaps_CP_641_symbol <= initIfMaps_CP_641_elements(233);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	78 
    -- CP-element group 0: 	79 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	149 
    -- CP-element group 0: 	152 
    -- CP-element group 0: 	133 
    -- CP-element group 0: 	134 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	127 
    -- CP-element group 0: 	128 
    -- CP-element group 0: 	131 
    -- CP-element group 0: 	123 
    -- CP-element group 0: 	165 
    -- CP-element group 0: 	167 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	96 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	139 
    -- CP-element group 0: 	180 
    -- CP-element group 0: 	181 
    -- CP-element group 0: 	183 
    -- CP-element group 0: 	124 
    -- CP-element group 0: 	126 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	87 
    -- CP-element group 0: 	88 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	118 
    -- CP-element group 0: 	120 
    -- CP-element group 0: 	102 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	159 
    -- CP-element group 0: 	160 
    -- CP-element group 0: 	162 
    -- CP-element group 0: 	136 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	141 
    -- CP-element group 0: 	142 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	178 
    -- CP-element group 0: 	99 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	94 
    -- CP-element group 0: 	111 
    -- CP-element group 0: 	112 
    -- CP-element group 0: 	146 
    -- CP-element group 0: 	147 
    -- CP-element group 0: 	170 
    -- CP-element group 0: 	108 
    -- CP-element group 0: 	168 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	157 
    -- CP-element group 0: 	173 
    -- CP-element group 0: 	172 
    -- CP-element group 0: 	90 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	106 
    -- CP-element group 0: 	154 
    -- CP-element group 0: 	155 
    -- CP-element group 0: 	114 
    -- CP-element group 0: 	144 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	175 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	42 
    -- CP-element group 0: 	43 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	54 
    -- CP-element group 0:  members (434) 
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Update/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Update/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Update/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Update/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_sample_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Sample/rr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Update/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Update/ccr
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_update_start_
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_resized_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_computed_1
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_259_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_268_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_272_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_281_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_285_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_294_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_223_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_536_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_380_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_211_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_223_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_509_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_355_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_491_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_399_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_217_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_217_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_374_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_437_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_520_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_495_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_502_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_502_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_255_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_351_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_412_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_418_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_482_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_446_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_370_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_552_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_229_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_229_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_235_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_235_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_389_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_450_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_568_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_456_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_393_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_431_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_469_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_465_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_361_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_427_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_478_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_408_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_211_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_298_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_304_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_313_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_317_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_323_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_332_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_336_store_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_342_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_259_store_0_req_1); -- 
    ccr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_268_call_req_1); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_272_store_0_req_1); -- 
    ccr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_281_call_req_1); -- 
    cr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_285_store_0_req_1); -- 
    ccr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_294_call_req_1); -- 
    rr_682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_223_inst_req_0); -- 
    ccr_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_536_call_req_1); -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_539_store_0_req_1); -- 
    req_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_539_index_offset_req_0); -- 
    req_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_512_index_offset_req_0); -- 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_512_index_offset_req_1); -- 
    cr_1256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_380_store_0_req_1); -- 
    rr_654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_211_inst_req_0); -- 
    cr_687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_223_inst_req_1); -- 
    ccr_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_509_call_req_1); -- 
    cr_1814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_512_store_0_req_1); -- 
    cr_1143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_355_store_0_req_1); -- 
    ccr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_491_call_req_1); -- 
    cr_1336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_399_store_0_req_1); -- 
    cr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_555_store_0_req_1); -- 
    req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_555_index_offset_req_0); -- 
    req_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_555_index_offset_req_1); -- 
    rr_668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_217_inst_req_0); -- 
    cr_673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_217_inst_req_1); -- 
    cr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_374_store_0_req_1); -- 
    cr_1496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_437_store_0_req_1); -- 
    cr_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_571_store_0_req_1); -- 
    req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_571_index_offset_req_0); -- 
    ccr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_520_call_req_1); -- 
    req_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_571_index_offset_req_1); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_495_store_0_req_1); -- 
    rr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_502_inst_req_0); -- 
    cr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_502_inst_req_1); -- 
    ccr_729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_255_call_req_1); -- 
    ccr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_351_call_req_1); -- 
    cr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_412_store_0_req_1); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_418_store_0_req_1); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_482_store_0_req_1); -- 
    ccr_1510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_446_call_req_1); -- 
    ccr_1190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_370_call_req_1); -- 
    req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_544_index_offset_req_1); -- 
    ccr_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_552_call_req_1); -- 
    cr_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_523_store_0_req_1); -- 
    req_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_523_index_offset_req_0); -- 
    rr_696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_229_inst_req_0); -- 
    cr_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_229_inst_req_1); -- 
    rr_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_235_inst_req_0); -- 
    cr_715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_235_inst_req_1); -- 
    req_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_523_index_offset_req_1); -- 
    ccr_1270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_389_call_req_1); -- 
    cr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_450_store_0_req_1); -- 
    ccr_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_568_call_req_1); -- 
    cr_1576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_456_store_0_req_1); -- 
    cr_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_393_store_0_req_1); -- 
    cr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_431_store_0_req_1); -- 
    cr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_469_store_0_req_1); -- 
    cr_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_560_store_0_req_1); -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_560_index_offset_req_0); -- 
    ccr_1590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_465_call_req_1); -- 
    cr_1176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_361_store_0_req_1); -- 
    cr_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_544_store_0_req_1); -- 
    req_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_544_index_offset_req_0); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_560_index_offset_req_1); -- 
    req_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_528_index_offset_req_0); -- 
    req_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_528_index_offset_req_1); -- 
    ccr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_427_call_req_1); -- 
    req_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_539_index_offset_req_1); -- 
    ccr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_478_call_req_1); -- 
    cr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_528_store_0_req_1); -- 
    ccr_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_408_call_req_1); -- 
    cr_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => type_cast_211_inst_req_1); -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_298_store_0_req_1); -- 
    cr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_304_store_0_req_1); -- 
    ccr_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_313_call_req_1); -- 
    cr_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_317_store_0_req_1); -- 
    cr_1016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_323_store_0_req_1); -- 
    ccr_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => call_stmt_332_call_req_1); -- 
    cr_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_336_store_0_req_1); -- 
    cr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(0), ack => array_obj_ref_342_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Sample/ra
      -- CP-element group 1: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_211_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_0, ack => initIfMaps_CP_641_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	129 
    -- CP-element group 2: 	11 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Update/ca
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_Update/$exit
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/type_cast_211_update_completed_
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Sample/crr
      -- CP-element group 2: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_211_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_255_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ca_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_211_inst_ack_1, ack => initIfMaps_CP_641_elements(2)); -- 
    crr_724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(2), ack => call_stmt_255_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Sample/ra
      -- CP-element group 3: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_217_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_217_inst_ack_0, ack => initIfMaps_CP_641_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	28 
    -- CP-element group 4: 	137 
    -- CP-element group 4: 	37 
    -- CP-element group 4: 	46 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Update/ca
      -- CP-element group 4: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_update_completed_
      -- CP-element group 4: 	 assign_stmt_208_to_assign_stmt_577/type_cast_217_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_217_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_217_inst_ack_1, ack => initIfMaps_CP_641_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Sample/ra
      -- CP-element group 5: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_223_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_223_inst_ack_0, ack => initIfMaps_CP_641_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	150 
    -- CP-element group 6: 	64 
    -- CP-element group 6: 	73 
    -- CP-element group 6: 	55 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Update/ca
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_Update/$exit
      -- CP-element group 6: 	 assign_stmt_208_to_assign_stmt_577/type_cast_223_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_223_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_223_inst_ack_1, ack => initIfMaps_CP_641_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Sample/ra
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_sample_completed_
      -- CP-element group 7: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_229_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_229_inst_ack_0, ack => initIfMaps_CP_641_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	100 
    -- CP-element group 8: 	163 
    -- CP-element group 8: 	91 
    -- CP-element group 8: 	82 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_update_completed_
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Update/$exit
      -- CP-element group 8: 	 assign_stmt_208_to_assign_stmt_577/type_cast_229_Update/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_229_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_229_inst_ack_1, ack => initIfMaps_CP_641_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_sample_completed_
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Sample/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_235_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_235_inst_ack_0, ack => initIfMaps_CP_641_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	121 
    -- CP-element group 10: 	176 
    -- CP-element group 10: 	109 
    -- CP-element group 10: 	115 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Update/ca
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_Update/$exit
      -- CP-element group 10: 	 assign_stmt_208_to_assign_stmt_577/type_cast_235_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_235_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_235_inst_ack_1, ack => initIfMaps_CP_641_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Sample/cra
      -- CP-element group 11: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_255_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_255_call_ack_0, ack => initIfMaps_CP_641_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	199 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Update/cca
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_update_completed_
      -- CP-element group 12: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_255_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_255_call_ack_1, ack => initIfMaps_CP_641_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_sample_start_
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/array_obj_ref_259_Split/$entry
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/array_obj_ref_259_Split/$exit
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/array_obj_ref_259_Split/split_req
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/array_obj_ref_259_Split/split_ack
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/$entry
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_259_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(13), ack => array_obj_ref_259_store_0_req_0); -- 
    initIfMaps_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(12) & initIfMaps_CP_641_elements(0);
      gj_initIfMaps_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	218 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_sample_completed_
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/$exit
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/$exit
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_259_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_259_store_0_ack_0, ack => initIfMaps_CP_641_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	233 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_update_completed_
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/$exit
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/$exit
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_259_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_259_store_0_ack_1, ack => initIfMaps_CP_641_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	199 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_sample_start_
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_268_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(16), ack => call_stmt_268_call_req_0); -- 
    initIfMaps_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(199) & initIfMaps_CP_641_elements(2);
      gj_initIfMaps_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_sample_completed_
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Sample/$exit
      -- CP-element group 17: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_268_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_268_call_ack_0, ack => initIfMaps_CP_641_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	200 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_update_completed_
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Update/$exit
      -- CP-element group 18: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_268_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_268_call_ack_1, ack => initIfMaps_CP_641_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	0 
    -- CP-element group 19: 	218 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_sample_start_
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/$entry
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/array_obj_ref_272_Split/$entry
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/array_obj_ref_272_Split/$exit
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/array_obj_ref_272_Split/split_req
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/array_obj_ref_272_Split/split_ack
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/$entry
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_272_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(19), ack => array_obj_ref_272_store_0_req_0); -- 
    initIfMaps_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(18) & initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(218);
      gj_initIfMaps_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	219 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_sample_completed_
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/$exit
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/$exit
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_272_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_272_store_0_ack_0, ack => initIfMaps_CP_641_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	233 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_update_completed_
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/$exit
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/$exit
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_272_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_272_store_0_ack_1, ack => initIfMaps_CP_641_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	200 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_sample_start_
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_281_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(22), ack => call_stmt_281_call_req_0); -- 
    initIfMaps_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(200) & initIfMaps_CP_641_elements(2);
      gj_initIfMaps_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_sample_completed_
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_281_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_281_call_ack_0, ack => initIfMaps_CP_641_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	201 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_update_completed_
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Update/$exit
      -- CP-element group 24: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_281_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_281_call_ack_1, ack => initIfMaps_CP_641_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: 	0 
    -- CP-element group 25: 	219 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_sample_start_
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/array_obj_ref_285_Split/$entry
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/array_obj_ref_285_Split/$exit
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/array_obj_ref_285_Split/split_req
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/array_obj_ref_285_Split/split_ack
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/$entry
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/word_0/$entry
      -- CP-element group 25: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_285_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(25), ack => array_obj_ref_285_store_0_req_0); -- 
    initIfMaps_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(24) & initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(219);
      gj_initIfMaps_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	220 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_sample_completed_
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/$exit
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/$exit
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/word_0/$exit
      -- CP-element group 26: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_285_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_285_store_0_ack_0, ack => initIfMaps_CP_641_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	233 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_update_completed_
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/$exit
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/$exit
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/word_0/$exit
      -- CP-element group 27: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_285_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_285_store_0_ack_1, ack => initIfMaps_CP_641_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	4 
    -- CP-element group 28: 	201 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_sample_start_
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Sample/$entry
      -- CP-element group 28: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_294_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(28), ack => call_stmt_294_call_req_0); -- 
    initIfMaps_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(4) & initIfMaps_CP_641_elements(201);
      gj_initIfMaps_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_sample_completed_
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_294_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_294_call_ack_0, ack => initIfMaps_CP_641_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	202 
    -- CP-element group 30: 	34 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_update_completed_
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Update/$exit
      -- CP-element group 30: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_294_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_294_call_ack_1, ack => initIfMaps_CP_641_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	0 
    -- CP-element group 31: 	220 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_sample_start_
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/$entry
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/array_obj_ref_298_Split/$entry
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/array_obj_ref_298_Split/$exit
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/array_obj_ref_298_Split/split_req
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/array_obj_ref_298_Split/split_ack
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/$entry
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_298_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(31), ack => array_obj_ref_298_store_0_req_0); -- 
    initIfMaps_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(30) & initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(220);
      gj_initIfMaps_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	221 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_sample_completed_
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/$exit
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_298_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_298_store_0_ack_0, ack => initIfMaps_CP_641_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	233 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_update_completed_
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/$exit
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/$exit
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_298_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_298_store_0_ack_1, ack => initIfMaps_CP_641_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	30 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_sample_start_
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/array_obj_ref_304_Split/$entry
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/array_obj_ref_304_Split/$exit
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/array_obj_ref_304_Split/split_req
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/array_obj_ref_304_Split/split_ack
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/$entry
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_304_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(34), ack => array_obj_ref_304_store_0_req_0); -- 
    initIfMaps_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(30) & initIfMaps_CP_641_elements(0);
      gj_initIfMaps_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	184 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_sample_completed_
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/$exit
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_304_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_0, ack => initIfMaps_CP_641_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	233 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_update_completed_
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/$exit
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/$exit
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_304_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_1, ack => initIfMaps_CP_641_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	4 
    -- CP-element group 37: 	202 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_sample_start_
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Sample/$entry
      -- CP-element group 37: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_313_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(37), ack => call_stmt_313_call_req_0); -- 
    initIfMaps_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(4) & initIfMaps_CP_641_elements(202);
      gj_initIfMaps_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_sample_completed_
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_313_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_313_call_ack_0, ack => initIfMaps_CP_641_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	203 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	43 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_update_completed_
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Update/$exit
      -- CP-element group 39: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_313_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_313_call_ack_1, ack => initIfMaps_CP_641_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: 	221 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_sample_start_
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/array_obj_ref_317_Split/$entry
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/array_obj_ref_317_Split/$exit
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/array_obj_ref_317_Split/split_req
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/array_obj_ref_317_Split/split_ack
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_317_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(40), ack => array_obj_ref_317_store_0_req_0); -- 
    initIfMaps_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(221) & initIfMaps_CP_641_elements(39);
      gj_initIfMaps_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	222 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_sample_completed_
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/$exit
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/$exit
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/word_0/$exit
      -- CP-element group 41: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_317_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_317_store_0_ack_0, ack => initIfMaps_CP_641_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	0 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	233 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_update_completed_
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/$exit
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/$exit
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_317_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_317_store_0_ack_1, ack => initIfMaps_CP_641_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	0 
    -- CP-element group 43: 	184 
    -- CP-element group 43: 	39 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_sample_start_
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/$entry
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/array_obj_ref_323_Split/$entry
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/array_obj_ref_323_Split/$exit
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/array_obj_ref_323_Split/split_req
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/array_obj_ref_323_Split/split_ack
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/$entry
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/word_0/$entry
      -- CP-element group 43: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_323_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(43), ack => array_obj_ref_323_store_0_req_0); -- 
    initIfMaps_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(184) & initIfMaps_CP_641_elements(39);
      gj_initIfMaps_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	185 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_sample_completed_
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/$exit
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/word_0/$exit
      -- CP-element group 44: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_323_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_323_store_0_ack_0, ack => initIfMaps_CP_641_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	233 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_update_completed_
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/$exit
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/$exit
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/word_0/$exit
      -- CP-element group 45: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_323_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_323_store_0_ack_1, ack => initIfMaps_CP_641_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	4 
    -- CP-element group 46: 	203 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_sample_start_
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Sample/$entry
      -- CP-element group 46: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_332_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(46), ack => call_stmt_332_call_req_0); -- 
    initIfMaps_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(4) & initIfMaps_CP_641_elements(203);
      gj_initIfMaps_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_sample_completed_
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Sample/$exit
      -- CP-element group 47: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_332_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_332_call_ack_0, ack => initIfMaps_CP_641_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	204 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	52 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_update_completed_
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Update/$exit
      -- CP-element group 48: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_332_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_332_call_ack_1, ack => initIfMaps_CP_641_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: 	222 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_sample_start_
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/$entry
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/array_obj_ref_336_Split/$entry
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/array_obj_ref_336_Split/$exit
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/array_obj_ref_336_Split/split_req
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/array_obj_ref_336_Split/split_ack
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/$entry
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_336_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(49), ack => array_obj_ref_336_store_0_req_0); -- 
    initIfMaps_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(222) & initIfMaps_CP_641_elements(48);
      gj_initIfMaps_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	223 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_sample_completed_
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_336_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_336_store_0_ack_0, ack => initIfMaps_CP_641_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	233 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_update_completed_
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/$exit
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_336_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_336_store_0_ack_1, ack => initIfMaps_CP_641_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: 	185 
    -- CP-element group 52: 	48 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_sample_start_
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/array_obj_ref_342_Split/$entry
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/array_obj_ref_342_Split/$exit
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/array_obj_ref_342_Split/split_req
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/array_obj_ref_342_Split/split_ack
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/$entry
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/word_0/$entry
      -- CP-element group 52: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_342_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(52), ack => array_obj_ref_342_store_0_req_0); -- 
    initIfMaps_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(185) & initIfMaps_CP_641_elements(48);
      gj_initIfMaps_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	186 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_sample_completed_
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/$exit
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/$exit
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/word_0/$exit
      -- CP-element group 53: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_342_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_342_store_0_ack_0, ack => initIfMaps_CP_641_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	233 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_update_completed_
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/$exit
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/$exit
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/word_0/$exit
      -- CP-element group 54: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_342_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_342_store_0_ack_1, ack => initIfMaps_CP_641_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	6 
    -- CP-element group 55: 	204 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_sample_start_
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Sample/$entry
      -- CP-element group 55: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_351_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(55), ack => call_stmt_351_call_req_0); -- 
    initIfMaps_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(6) & initIfMaps_CP_641_elements(204);
      gj_initIfMaps_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_sample_completed_
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Sample/$exit
      -- CP-element group 56: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_351_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_351_call_ack_0, ack => initIfMaps_CP_641_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	205 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_update_completed_
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Update/$exit
      -- CP-element group 57: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_351_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_351_call_ack_1, ack => initIfMaps_CP_641_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	223 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_sample_start_
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/$entry
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/array_obj_ref_355_Split/$entry
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/array_obj_ref_355_Split/$exit
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/array_obj_ref_355_Split/split_req
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/array_obj_ref_355_Split/split_ack
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/$entry
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_355_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(58), ack => array_obj_ref_355_store_0_req_0); -- 
    initIfMaps_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(57) & initIfMaps_CP_641_elements(223);
      gj_initIfMaps_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	224 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_sample_completed_
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/$exit
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/$exit
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_355_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_355_store_0_ack_0, ack => initIfMaps_CP_641_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	233 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_update_completed_
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/$exit
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/$exit
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_355_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_355_store_0_ack_1, ack => initIfMaps_CP_641_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: 	57 
    -- CP-element group 61: 	186 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_sample_start_
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/$entry
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/array_obj_ref_361_Split/$entry
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/array_obj_ref_361_Split/$exit
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/array_obj_ref_361_Split/split_req
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/array_obj_ref_361_Split/split_ack
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/$entry
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_361_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(61), ack => array_obj_ref_361_store_0_req_0); -- 
    initIfMaps_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(57) & initIfMaps_CP_641_elements(186);
      gj_initIfMaps_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	187 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_sample_completed_
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/$exit
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_361_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_361_store_0_ack_0, ack => initIfMaps_CP_641_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	233 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_update_completed_
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/$exit
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/$exit
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_361_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_361_store_0_ack_1, ack => initIfMaps_CP_641_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	6 
    -- CP-element group 64: 	205 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_sample_start_
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_370_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(64), ack => call_stmt_370_call_req_0); -- 
    initIfMaps_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(6) & initIfMaps_CP_641_elements(205);
      gj_initIfMaps_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_sample_completed_
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Sample/$exit
      -- CP-element group 65: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_370_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_370_call_ack_0, ack => initIfMaps_CP_641_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	70 
    -- CP-element group 66: 	206 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_update_completed_
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Update/$exit
      -- CP-element group 66: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_370_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_370_call_ack_1, ack => initIfMaps_CP_641_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: 	66 
    -- CP-element group 67: 	224 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_sample_start_
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/$entry
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/array_obj_ref_374_Split/$entry
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/array_obj_ref_374_Split/$exit
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/array_obj_ref_374_Split/split_req
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/array_obj_ref_374_Split/split_ack
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/$entry
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/word_0/$entry
      -- CP-element group 67: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_374_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(67), ack => array_obj_ref_374_store_0_req_0); -- 
    initIfMaps_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(66) & initIfMaps_CP_641_elements(224);
      gj_initIfMaps_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	225 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_sample_completed_
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/$exit
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/$exit
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/word_0/$exit
      -- CP-element group 68: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_374_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_374_store_0_ack_0, ack => initIfMaps_CP_641_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	233 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_update_completed_
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/$exit
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/$exit
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_374_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_374_store_0_ack_1, ack => initIfMaps_CP_641_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: 	66 
    -- CP-element group 70: 	187 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_sample_start_
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/$entry
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/array_obj_ref_380_Split/$entry
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/array_obj_ref_380_Split/$exit
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/array_obj_ref_380_Split/split_req
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/array_obj_ref_380_Split/split_ack
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/$entry
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/word_0/$entry
      -- CP-element group 70: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_380_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(70), ack => array_obj_ref_380_store_0_req_0); -- 
    initIfMaps_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(66) & initIfMaps_CP_641_elements(187);
      gj_initIfMaps_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	188 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_sample_completed_
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/$exit
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/$exit
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/word_0/$exit
      -- CP-element group 71: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_380_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_380_store_0_ack_0, ack => initIfMaps_CP_641_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	233 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_update_completed_
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/$exit
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/$exit
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/word_0/$exit
      -- CP-element group 72: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_380_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_380_store_0_ack_1, ack => initIfMaps_CP_641_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	6 
    -- CP-element group 73: 	206 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_sample_start_
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Sample/$entry
      -- CP-element group 73: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_389_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(73), ack => call_stmt_389_call_req_0); -- 
    initIfMaps_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(6) & initIfMaps_CP_641_elements(206);
      gj_initIfMaps_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_sample_completed_
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_389_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_389_call_ack_0, ack => initIfMaps_CP_641_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	207 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_update_completed_
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Update/$exit
      -- CP-element group 75: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_389_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_389_call_ack_1, ack => initIfMaps_CP_641_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: 	225 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/word_0/rr
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/word_0/$entry
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_sample_start_
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/array_obj_ref_393_Split/$entry
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/array_obj_ref_393_Split/$exit
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/array_obj_ref_393_Split/split_req
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/array_obj_ref_393_Split/split_ack
      -- CP-element group 76: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_393_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(76), ack => array_obj_ref_393_store_0_req_0); -- 
    initIfMaps_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(225) & initIfMaps_CP_641_elements(75);
      gj_initIfMaps_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	226 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/word_0/ra
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/word_0/$exit
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_sample_completed_
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/$exit
      -- CP-element group 77: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_393_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_393_store_0_ack_0, ack => initIfMaps_CP_641_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	0 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	233 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/word_0/$exit
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/word_0/ca
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/$exit
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_Update/word_access_complete/$exit
      -- CP-element group 78: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_393_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_393_store_0_ack_1, ack => initIfMaps_CP_641_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	0 
    -- CP-element group 79: 	188 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/word_0/rr
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_sample_start_
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/word_0/$entry
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/$entry
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/array_obj_ref_399_Split/$exit
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/array_obj_ref_399_Split/$entry
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/$entry
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/array_obj_ref_399_Split/split_req
      -- CP-element group 79: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/array_obj_ref_399_Split/split_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_399_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(79), ack => array_obj_ref_399_store_0_req_0); -- 
    initIfMaps_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(188) & initIfMaps_CP_641_elements(75);
      gj_initIfMaps_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	189 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/$exit
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_sample_completed_
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/word_0/$exit
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/word_0/ra
      -- CP-element group 80: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_399_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_399_store_0_ack_0, ack => initIfMaps_CP_641_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	233 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/$exit
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/word_0/ca
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/$exit
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_Update/word_access_complete/word_0/$exit
      -- CP-element group 81: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_399_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_399_store_0_ack_1, ack => initIfMaps_CP_641_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	207 
    -- CP-element group 82: 	8 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Sample/crr
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Sample/$entry
      -- CP-element group 82: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_408_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(82), ack => call_stmt_408_call_req_0); -- 
    initIfMaps_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(207) & initIfMaps_CP_641_elements(8);
      gj_initIfMaps_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_sample_completed_
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Sample/$exit
      -- CP-element group 83: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_408_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_408_call_ack_0, ack => initIfMaps_CP_641_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	208 
    -- CP-element group 84: 	88 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_update_completed_
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Update/$exit
      -- CP-element group 84: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_408_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_408_call_ack_1, ack => initIfMaps_CP_641_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: 	226 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/word_0/rr
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/word_0/$entry
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/$entry
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/array_obj_ref_412_Split/split_ack
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/array_obj_ref_412_Split/split_req
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/array_obj_ref_412_Split/$exit
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/array_obj_ref_412_Split/$entry
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/$entry
      -- CP-element group 85: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_412_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(85), ack => array_obj_ref_412_store_0_req_0); -- 
    initIfMaps_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(226) & initIfMaps_CP_641_elements(84);
      gj_initIfMaps_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	227 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/word_0/ra
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/word_0/$exit
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/word_access_start/$exit
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_412_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_412_store_0_ack_0, ack => initIfMaps_CP_641_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	0 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	233 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/word_0/ca
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/word_0/$exit
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/word_access_complete/$exit
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_Update/$exit
      -- CP-element group 87: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_412_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_412_store_0_ack_1, ack => initIfMaps_CP_641_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	0 
    -- CP-element group 88: 	189 
    -- CP-element group 88: 	84 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/word_0/rr
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/word_0/$entry
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/$entry
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/array_obj_ref_418_Split/split_ack
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/array_obj_ref_418_Split/split_req
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/array_obj_ref_418_Split/$exit
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/array_obj_ref_418_Split/$entry
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_418_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(88), ack => array_obj_ref_418_store_0_req_0); -- 
    initIfMaps_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(189) & initIfMaps_CP_641_elements(84);
      gj_initIfMaps_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	190 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/word_0/ra
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/word_0/$exit
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/word_access_start/$exit
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Sample/$exit
      -- CP-element group 89: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_418_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_418_store_0_ack_0, ack => initIfMaps_CP_641_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	0 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	233 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/word_0/ca
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/word_0/$exit
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/word_access_complete/$exit
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_Update/$exit
      -- CP-element group 90: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_418_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_418_store_0_ack_1, ack => initIfMaps_CP_641_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	208 
    -- CP-element group 91: 	8 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Sample/$entry
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Sample/crr
      -- CP-element group 91: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_427_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(91), ack => call_stmt_427_call_req_0); -- 
    initIfMaps_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(208) & initIfMaps_CP_641_elements(8);
      gj_initIfMaps_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Sample/cra
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Sample/$exit
      -- CP-element group 92: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_427_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_427_call_ack_0, ack => initIfMaps_CP_641_elements(92)); -- 
    -- CP-element group 93:  fork  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	209 
    -- CP-element group 93: 	97 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Update/cca
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_update_completed_
      -- CP-element group 93: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_427_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_427_call_ack_1, ack => initIfMaps_CP_641_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	0 
    -- CP-element group 94: 	227 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/$entry
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/$entry
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/array_obj_ref_431_Split/split_req
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/array_obj_ref_431_Split/split_ack
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/array_obj_ref_431_Split/$exit
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_sample_start_
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/array_obj_ref_431_Split/$entry
      -- CP-element group 94: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_431_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(94), ack => array_obj_ref_431_store_0_req_0); -- 
    initIfMaps_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(227) & initIfMaps_CP_641_elements(93);
      gj_initIfMaps_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	228 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/$exit
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/$exit
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_sample_completed_
      -- CP-element group 95: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_431_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_431_store_0_ack_0, ack => initIfMaps_CP_641_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	0 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	233 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_update_completed_
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/word_access_complete/$exit
      -- CP-element group 96: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_431_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_431_store_0_ack_1, ack => initIfMaps_CP_641_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: 	190 
    -- CP-element group 97: 	93 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/array_obj_ref_437_Split/split_req
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/array_obj_ref_437_Split/$entry
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/$entry
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/array_obj_ref_437_Split/$exit
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/$entry
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_sample_start_
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/word_0/rr
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/array_obj_ref_437_Split/split_ack
      -- CP-element group 97: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/word_0/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_437_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(97), ack => array_obj_ref_437_store_0_req_0); -- 
    initIfMaps_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "initIfMaps_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(190) & initIfMaps_CP_641_elements(93);
      gj_initIfMaps_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	191 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/word_0/ra
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/$exit
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_sample_completed_
      -- CP-element group 98: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_437_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_437_store_0_ack_0, ack => initIfMaps_CP_641_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	0 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	233 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_update_completed_
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/$exit
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/word_0/$exit
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/$exit
      -- CP-element group 99: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_437_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_437_store_0_ack_1, ack => initIfMaps_CP_641_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	209 
    -- CP-element group 100: 	8 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Sample/crr
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_sample_start_
      -- CP-element group 100: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Sample/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_446_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(100), ack => call_stmt_446_call_req_0); -- 
    initIfMaps_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(209) & initIfMaps_CP_641_elements(8);
      gj_initIfMaps_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Sample/cra
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_sample_completed_
      -- CP-element group 101: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_446_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_446_call_ack_0, ack => initIfMaps_CP_641_elements(101)); -- 
    -- CP-element group 102:  fork  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	0 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	210 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	106 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Update/cca
      -- CP-element group 102: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_update_completed_
      -- CP-element group 102: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_446_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_446_call_ack_1, ack => initIfMaps_CP_641_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: 	228 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/word_0/$entry
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/word_0/rr
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/array_obj_ref_450_Split/split_ack
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_sample_start_
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/$entry
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/array_obj_ref_450_Split/split_req
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/$entry
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/array_obj_ref_450_Split/$exit
      -- CP-element group 103: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/array_obj_ref_450_Split/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_450_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(103), ack => array_obj_ref_450_store_0_req_0); -- 
    initIfMaps_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(228) & initIfMaps_CP_641_elements(102);
      gj_initIfMaps_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	229 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_sample_completed_
      -- CP-element group 104: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/$exit
      -- CP-element group 104: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/word_0/$exit
      -- CP-element group 104: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/word_access_start/word_0/ra
      -- CP-element group 104: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_450_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_store_0_ack_0, ack => initIfMaps_CP_641_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	233 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/word_0/$exit
      -- CP-element group 105: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_update_completed_
      -- CP-element group 105: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/word_0/ca
      -- CP-element group 105: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/word_access_complete/$exit
      -- CP-element group 105: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_450_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_450_store_0_ack_1, ack => initIfMaps_CP_641_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	0 
    -- CP-element group 106: 	191 
    -- CP-element group 106: 	102 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/array_obj_ref_456_Split/split_req
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/array_obj_ref_456_Split/split_ack
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/$entry
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/array_obj_ref_456_Split/$exit
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_sample_start_
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/$entry
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/word_0/$entry
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/array_obj_ref_456_Split/$entry
      -- CP-element group 106: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_456_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(106), ack => array_obj_ref_456_store_0_req_0); -- 
    initIfMaps_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(191) & initIfMaps_CP_641_elements(102);
      gj_initIfMaps_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	192 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/$exit
      -- CP-element group 107: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/$exit
      -- CP-element group 107: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/word_0/ra
      -- CP-element group 107: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_sample_completed_
      -- CP-element group 107: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_456_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_456_store_0_ack_0, ack => initIfMaps_CP_641_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	0 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	233 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_update_completed_
      -- CP-element group 108: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/$exit
      -- CP-element group 108: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/$exit
      -- CP-element group 108: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_456_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_456_store_0_ack_1, ack => initIfMaps_CP_641_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	210 
    -- CP-element group 109: 	10 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Sample/crr
      -- CP-element group 109: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_sample_start_
      -- CP-element group 109: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Sample/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_465_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(109), ack => call_stmt_465_call_req_0); -- 
    initIfMaps_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(210) & initIfMaps_CP_641_elements(10);
      gj_initIfMaps_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Sample/cra
      -- CP-element group 110: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_sample_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_465_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_465_call_ack_0, ack => initIfMaps_CP_641_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	0 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	211 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Update/cca
      -- CP-element group 111: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_Update/$exit
      -- CP-element group 111: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_465_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_465_call_ack_1, ack => initIfMaps_CP_641_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	0 
    -- CP-element group 112: 	192 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/word_0/$entry
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/word_0/rr
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/array_obj_ref_469_Split/split_ack
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_sample_start_
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/$entry
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/array_obj_ref_469_Split/split_req
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/array_obj_ref_469_Split/$entry
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/array_obj_ref_469_Split/$exit
      -- CP-element group 112: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_469_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(112), ack => array_obj_ref_469_store_0_req_0); -- 
    initIfMaps_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(192) & initIfMaps_CP_641_elements(111);
      gj_initIfMaps_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	193 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/word_0/$exit
      -- CP-element group 113: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/word_0/ra
      -- CP-element group 113: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_sample_completed_
      -- CP-element group 113: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/word_access_start/$exit
      -- CP-element group 113: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_469_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_469_store_0_ack_0, ack => initIfMaps_CP_641_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	0 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	233 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_update_completed_
      -- CP-element group 114: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/$exit
      -- CP-element group 114: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/$exit
      -- CP-element group 114: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_469_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_469_store_0_ack_1, ack => initIfMaps_CP_641_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	211 
    -- CP-element group 115: 	10 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_sample_start_
      -- CP-element group 115: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Sample/crr
      -- CP-element group 115: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Sample/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_478_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(115), ack => call_stmt_478_call_req_0); -- 
    initIfMaps_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(211) & initIfMaps_CP_641_elements(10);
      gj_initIfMaps_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_sample_completed_
      -- CP-element group 116: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Sample/cra
      -- CP-element group 116: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_478_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_478_call_ack_0, ack => initIfMaps_CP_641_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	212 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Update/cca
      -- CP-element group 117: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_update_completed_
      -- CP-element group 117: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_Update/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_478_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_478_call_ack_1, ack => initIfMaps_CP_641_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	0 
    -- CP-element group 118: 	193 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/array_obj_ref_482_Split/split_req
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/array_obj_ref_482_Split/split_ack
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/word_0/rr
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/$entry
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_sample_start_
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/$entry
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/array_obj_ref_482_Split/$entry
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/array_obj_ref_482_Split/$exit
      -- CP-element group 118: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/word_0/$entry
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_482_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(118), ack => array_obj_ref_482_store_0_req_0); -- 
    initIfMaps_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(193) & initIfMaps_CP_641_elements(117);
      gj_initIfMaps_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	194 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/word_0/ra
      -- CP-element group 119: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_sample_completed_
      -- CP-element group 119: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/$exit
      -- CP-element group 119: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_482_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_store_0_ack_0, ack => initIfMaps_CP_641_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	0 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	233 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/$exit
      -- CP-element group 120: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_Update/word_access_complete/$exit
      -- CP-element group 120: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_482_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_482_store_0_ack_1, ack => initIfMaps_CP_641_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	212 
    -- CP-element group 121: 	10 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Sample/crr
      -- CP-element group 121: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Sample/$entry
      -- CP-element group 121: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_sample_start_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_491_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(121), ack => call_stmt_491_call_req_0); -- 
    initIfMaps_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(212) & initIfMaps_CP_641_elements(10);
      gj_initIfMaps_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Sample/cra
      -- CP-element group 122: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_sample_completed_
      -- CP-element group 122: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Sample/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_491_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_491_call_ack_0, ack => initIfMaps_CP_641_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	0 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	213 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Update/$exit
      -- CP-element group 123: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_Update/cca
      -- CP-element group 123: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_update_completed_
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_491_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_491_call_ack_1, ack => initIfMaps_CP_641_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	0 
    -- CP-element group 124: 	194 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/array_obj_ref_495_Split/$exit
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_sample_start_
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/word_0/$entry
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/array_obj_ref_495_Split/split_req
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/array_obj_ref_495_Split/$entry
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/$entry
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/array_obj_ref_495_Split/split_ack
      -- CP-element group 124: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_495_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(124), ack => array_obj_ref_495_store_0_req_0); -- 
    initIfMaps_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(0) & initIfMaps_CP_641_elements(194) & initIfMaps_CP_641_elements(123);
      gj_initIfMaps_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	195 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_sample_completed_
      -- CP-element group 125: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/word_0/ra
      -- CP-element group 125: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/$exit
      -- CP-element group 125: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_495_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_495_store_0_ack_0, ack => initIfMaps_CP_641_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	0 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	233 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_update_completed_
      -- CP-element group 126: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/$exit
      -- CP-element group 126: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/$exit
      -- CP-element group 126: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_495_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_495_store_0_ack_1, ack => initIfMaps_CP_641_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	0 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_sample_completed_
      -- CP-element group 127: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Sample/$exit
      -- CP-element group 127: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Sample/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_502_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_0, ack => initIfMaps_CP_641_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	0 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	150 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	137 
    -- CP-element group 128: 	163 
    -- CP-element group 128: 	176 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_update_completed_
      -- CP-element group 128: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Update/$exit
      -- CP-element group 128: 	 assign_stmt_208_to_assign_stmt_577/type_cast_502_Update/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:type_cast_502_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_1, ack => initIfMaps_CP_641_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	213 
    -- CP-element group 129: 	2 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_sample_start_
      -- CP-element group 129: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Sample/$entry
      -- CP-element group 129: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_509_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(129), ack => call_stmt_509_call_req_0); -- 
    initIfMaps_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(128) & initIfMaps_CP_641_elements(213) & initIfMaps_CP_641_elements(2);
      gj_initIfMaps_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_sample_completed_
      -- CP-element group 130: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Sample/$exit
      -- CP-element group 130: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_509_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_509_call_ack_0, ack => initIfMaps_CP_641_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	0 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	214 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_update_completed_
      -- CP-element group 131: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Update/$exit
      -- CP-element group 131: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_509_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_509_call_ack_1, ack => initIfMaps_CP_641_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: 	131 
    -- CP-element group 132: 	229 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	135 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_sample_start_
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/$entry
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/array_obj_ref_512_Split/$entry
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/array_obj_ref_512_Split/$exit
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/array_obj_ref_512_Split/split_req
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/array_obj_ref_512_Split/split_ack
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/$entry
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/word_0/$entry
      -- CP-element group 132: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(132), ack => array_obj_ref_512_store_0_req_0); -- 
    initIfMaps_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(134) & initIfMaps_CP_641_elements(131) & initIfMaps_CP_641_elements(229);
      gj_initIfMaps_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	0 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	233 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_sample_complete
      -- CP-element group 133: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Sample/$exit
      -- CP-element group 133: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_512_index_offset_ack_0, ack => initIfMaps_CP_641_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	0 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (13) 
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_word_address_calculated
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_root_address_calculated
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_offset_calculated
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Update/$exit
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_final_index_sum_regn_Update/ack
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_base_plus_offset/$entry
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_base_plus_offset/$exit
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_word_addrgen/$entry
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_word_addrgen/$exit
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_word_addrgen/root_register_req
      -- CP-element group 134: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_512_index_offset_ack_1, ack => initIfMaps_CP_641_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	132 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	230 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_sample_completed_
      -- CP-element group 135: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/$exit
      -- CP-element group 135: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/$exit
      -- CP-element group 135: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/word_0/$exit
      -- CP-element group 135: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_512_store_0_ack_0, ack => initIfMaps_CP_641_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	0 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	233 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_update_completed_
      -- CP-element group 136: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/$exit
      -- CP-element group 136: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/$exit
      -- CP-element group 136: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/word_0/$exit
      -- CP-element group 136: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_512_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_512_store_0_ack_1, ack => initIfMaps_CP_641_elements(136)); -- 
    -- CP-element group 137:  join  transition  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	4 
    -- CP-element group 137: 	128 
    -- CP-element group 137: 	214 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_sample_start_
      -- CP-element group 137: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Sample/$entry
      -- CP-element group 137: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_520_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(137), ack => call_stmt_520_call_req_0); -- 
    initIfMaps_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(4) & initIfMaps_CP_641_elements(128) & initIfMaps_CP_641_elements(214);
      gj_initIfMaps_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_sample_completed_
      -- CP-element group 138: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_520_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_520_call_ack_0, ack => initIfMaps_CP_641_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	0 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	215 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	145 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_update_completed_
      -- CP-element group 139: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Update/$exit
      -- CP-element group 139: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_520_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_520_call_ack_1, ack => initIfMaps_CP_641_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: 	230 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	143 
    -- CP-element group 140:  members (9) 
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_sample_start_
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/$entry
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/array_obj_ref_523_Split/$entry
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/array_obj_ref_523_Split/$exit
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/array_obj_ref_523_Split/split_req
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/array_obj_ref_523_Split/split_ack
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/$entry
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/word_0/$entry
      -- CP-element group 140: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(140), ack => array_obj_ref_523_store_0_req_0); -- 
    initIfMaps_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(139) & initIfMaps_CP_641_elements(230) & initIfMaps_CP_641_elements(142);
      gj_initIfMaps_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	0 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	233 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_sample_complete
      -- CP-element group 141: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Sample/$exit
      -- CP-element group 141: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_523_index_offset_ack_0, ack => initIfMaps_CP_641_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	0 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (13) 
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_word_address_calculated
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_root_address_calculated
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_offset_calculated
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Update/$exit
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_final_index_sum_regn_Update/ack
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_base_plus_offset/$entry
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_base_plus_offset/$exit
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_word_addrgen/$entry
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_word_addrgen/$exit
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_word_addrgen/root_register_req
      -- CP-element group 142: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_523_index_offset_ack_1, ack => initIfMaps_CP_641_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	140 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	231 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_sample_completed_
      -- CP-element group 143: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/$exit
      -- CP-element group 143: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/$exit
      -- CP-element group 143: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/word_0/$exit
      -- CP-element group 143: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_523_store_0_ack_0, ack => initIfMaps_CP_641_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	0 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	233 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_update_completed_
      -- CP-element group 144: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/$exit
      -- CP-element group 144: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/$exit
      -- CP-element group 144: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/word_0/$exit
      -- CP-element group 144: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_523_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_523_store_0_ack_1, ack => initIfMaps_CP_641_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	195 
    -- CP-element group 145: 	139 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	148 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_sample_start_
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/$entry
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/array_obj_ref_528_Split/$entry
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/array_obj_ref_528_Split/$exit
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/array_obj_ref_528_Split/split_req
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/array_obj_ref_528_Split/split_ack
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/$entry
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/word_0/$entry
      -- CP-element group 145: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(145), ack => array_obj_ref_528_store_0_req_0); -- 
    initIfMaps_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(195) & initIfMaps_CP_641_elements(139) & initIfMaps_CP_641_elements(147);
      gj_initIfMaps_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	0 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	233 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_sample_complete
      -- CP-element group 146: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Sample/$exit
      -- CP-element group 146: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_index_offset_ack_0, ack => initIfMaps_CP_641_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	0 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (13) 
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_word_address_calculated
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_root_address_calculated
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_offset_calculated
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Update/$exit
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_final_index_sum_regn_Update/ack
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_base_plus_offset/$entry
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_base_plus_offset/$exit
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_base_plus_offset/sum_rename_req
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_base_plus_offset/sum_rename_ack
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_word_addrgen/$entry
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_word_addrgen/$exit
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_word_addrgen/root_register_req
      -- CP-element group 147: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_index_offset_ack_1, ack => initIfMaps_CP_641_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	145 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	196 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_sample_completed_
      -- CP-element group 148: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/$exit
      -- CP-element group 148: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/$exit
      -- CP-element group 148: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/word_0/$exit
      -- CP-element group 148: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_store_0_ack_0, ack => initIfMaps_CP_641_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	0 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	233 
    -- CP-element group 149:  members (5) 
      -- CP-element group 149: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_update_completed_
      -- CP-element group 149: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/$exit
      -- CP-element group 149: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/$exit
      -- CP-element group 149: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/word_0/$exit
      -- CP-element group 149: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_528_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_528_store_0_ack_1, ack => initIfMaps_CP_641_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	6 
    -- CP-element group 150: 	128 
    -- CP-element group 150: 	215 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_sample_start_
      -- CP-element group 150: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Sample/$entry
      -- CP-element group 150: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_536_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(150), ack => call_stmt_536_call_req_0); -- 
    initIfMaps_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(6) & initIfMaps_CP_641_elements(128) & initIfMaps_CP_641_elements(215);
      gj_initIfMaps_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_sample_completed_
      -- CP-element group 151: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Sample/$exit
      -- CP-element group 151: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_536_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_536_call_ack_0, ack => initIfMaps_CP_641_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	0 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	216 
    -- CP-element group 152: 	158 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_update_completed_
      -- CP-element group 152: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Update/$exit
      -- CP-element group 152: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_536_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_536_call_ack_1, ack => initIfMaps_CP_641_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: 	231 
    -- CP-element group 153: 	155 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	156 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_sample_start_
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/$entry
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/array_obj_ref_539_Split/$entry
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/array_obj_ref_539_Split/$exit
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/array_obj_ref_539_Split/split_req
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/array_obj_ref_539_Split/split_ack
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/$entry
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/word_0/$entry
      -- CP-element group 153: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(153), ack => array_obj_ref_539_store_0_req_0); -- 
    initIfMaps_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(152) & initIfMaps_CP_641_elements(231) & initIfMaps_CP_641_elements(155);
      gj_initIfMaps_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	0 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	233 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_sample_complete
      -- CP-element group 154: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Sample/$exit
      -- CP-element group 154: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_index_offset_ack_0, ack => initIfMaps_CP_641_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	0 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (13) 
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_word_address_calculated
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_root_address_calculated
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_offset_calculated
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Update/$exit
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_final_index_sum_regn_Update/ack
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_base_plus_offset/$entry
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_base_plus_offset/$exit
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_base_plus_offset/sum_rename_req
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_base_plus_offset/sum_rename_ack
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_word_addrgen/$entry
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_word_addrgen/$exit
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_word_addrgen/root_register_req
      -- CP-element group 155: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_index_offset_ack_1, ack => initIfMaps_CP_641_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	232 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_sample_completed_
      -- CP-element group 156: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/$exit
      -- CP-element group 156: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/$exit
      -- CP-element group 156: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/word_0/$exit
      -- CP-element group 156: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_store_0_ack_0, ack => initIfMaps_CP_641_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	0 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	233 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_update_completed_
      -- CP-element group 157: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/$exit
      -- CP-element group 157: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/$exit
      -- CP-element group 157: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/word_0/$exit
      -- CP-element group 157: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_539_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_539_store_0_ack_1, ack => initIfMaps_CP_641_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	152 
    -- CP-element group 158: 	196 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	161 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_sample_start_
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/$entry
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/array_obj_ref_544_Split/$entry
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/array_obj_ref_544_Split/$exit
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/array_obj_ref_544_Split/split_req
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/array_obj_ref_544_Split/split_ack
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/$entry
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/word_0/$entry
      -- CP-element group 158: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(158), ack => array_obj_ref_544_store_0_req_0); -- 
    initIfMaps_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(152) & initIfMaps_CP_641_elements(196) & initIfMaps_CP_641_elements(160);
      gj_initIfMaps_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	0 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	233 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_sample_complete
      -- CP-element group 159: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Sample/$exit
      -- CP-element group 159: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_544_index_offset_ack_0, ack => initIfMaps_CP_641_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	0 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (13) 
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_word_address_calculated
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_root_address_calculated
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_offset_calculated
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Update/$exit
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_final_index_sum_regn_Update/ack
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_base_plus_offset/$entry
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_base_plus_offset/$exit
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_base_plus_offset/sum_rename_req
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_base_plus_offset/sum_rename_ack
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_word_addrgen/$entry
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_word_addrgen/$exit
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_word_addrgen/root_register_req
      -- CP-element group 160: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_544_index_offset_ack_1, ack => initIfMaps_CP_641_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	158 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	197 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_sample_completed_
      -- CP-element group 161: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/$exit
      -- CP-element group 161: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/$exit
      -- CP-element group 161: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/word_0/$exit
      -- CP-element group 161: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_544_store_0_ack_0, ack => initIfMaps_CP_641_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	0 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	233 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_update_completed_
      -- CP-element group 162: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/$exit
      -- CP-element group 162: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/$exit
      -- CP-element group 162: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/word_0/$exit
      -- CP-element group 162: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_544_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_544_store_0_ack_1, ack => initIfMaps_CP_641_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	128 
    -- CP-element group 163: 	216 
    -- CP-element group 163: 	8 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_sample_start_
      -- CP-element group 163: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Sample/$entry
      -- CP-element group 163: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_552_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(163), ack => call_stmt_552_call_req_0); -- 
    initIfMaps_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(128) & initIfMaps_CP_641_elements(216) & initIfMaps_CP_641_elements(8);
      gj_initIfMaps_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_sample_completed_
      -- CP-element group 164: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Sample/$exit
      -- CP-element group 164: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_552_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_552_call_ack_0, ack => initIfMaps_CP_641_elements(164)); -- 
    -- CP-element group 165:  fork  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	0 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	217 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	171 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_update_completed_
      -- CP-element group 165: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Update/$exit
      -- CP-element group 165: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_552_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_552_call_ack_1, ack => initIfMaps_CP_641_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: 	232 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	169 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_sample_start_
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/$entry
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/array_obj_ref_555_Split/$entry
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/array_obj_ref_555_Split/$exit
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/array_obj_ref_555_Split/split_req
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/array_obj_ref_555_Split/split_ack
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/$entry
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/word_0/$entry
      -- CP-element group 166: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(166), ack => array_obj_ref_555_store_0_req_0); -- 
    initIfMaps_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(165) & initIfMaps_CP_641_elements(232) & initIfMaps_CP_641_elements(168);
      gj_initIfMaps_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	0 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	233 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_sample_complete
      -- CP-element group 167: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_555_index_offset_ack_0, ack => initIfMaps_CP_641_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	0 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (13) 
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_word_address_calculated
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_root_address_calculated
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_offset_calculated
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_base_plus_offset/$entry
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_base_plus_offset/$exit
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_word_addrgen/$entry
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_word_addrgen/$exit
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_word_addrgen/root_register_req
      -- CP-element group 168: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_555_index_offset_ack_1, ack => initIfMaps_CP_641_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	166 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_sample_completed_
      -- CP-element group 169: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/$exit
      -- CP-element group 169: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/$exit
      -- CP-element group 169: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/word_0/$exit
      -- CP-element group 169: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_555_store_0_ack_0, ack => initIfMaps_CP_641_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	0 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	233 
    -- CP-element group 170:  members (5) 
      -- CP-element group 170: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_update_completed_
      -- CP-element group 170: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/$exit
      -- CP-element group 170: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/$exit
      -- CP-element group 170: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/word_0/$exit
      -- CP-element group 170: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_555_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_555_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_555_store_0_ack_1, ack => initIfMaps_CP_641_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	197 
    -- CP-element group 171: 	165 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	174 
    -- CP-element group 171:  members (9) 
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_sample_start_
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/$entry
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/array_obj_ref_560_Split/$entry
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/array_obj_ref_560_Split/$exit
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/array_obj_ref_560_Split/split_req
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/array_obj_ref_560_Split/split_ack
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/$entry
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/word_0/$entry
      -- CP-element group 171: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(171), ack => array_obj_ref_560_store_0_req_0); -- 
    initIfMaps_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(197) & initIfMaps_CP_641_elements(165) & initIfMaps_CP_641_elements(173);
      gj_initIfMaps_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	0 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	233 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_sample_complete
      -- CP-element group 172: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Sample/$exit
      -- CP-element group 172: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_560_index_offset_ack_0, ack => initIfMaps_CP_641_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	0 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (13) 
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_word_address_calculated
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_root_address_calculated
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_offset_calculated
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Update/$exit
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_final_index_sum_regn_Update/ack
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_base_plus_offset/$entry
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_base_plus_offset/$exit
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_word_addrgen/$entry
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_word_addrgen/$exit
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_word_addrgen/root_register_req
      -- CP-element group 173: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_560_index_offset_ack_1, ack => initIfMaps_CP_641_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	171 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	198 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_sample_completed_
      -- CP-element group 174: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/$exit
      -- CP-element group 174: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/$exit
      -- CP-element group 174: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/word_0/$exit
      -- CP-element group 174: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_560_store_0_ack_0, ack => initIfMaps_CP_641_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	0 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	233 
    -- CP-element group 175:  members (5) 
      -- CP-element group 175: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_update_completed_
      -- CP-element group 175: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/$exit
      -- CP-element group 175: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/$exit
      -- CP-element group 175: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/word_0/$exit
      -- CP-element group 175: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_560_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_560_store_0_ack_1, ack => initIfMaps_CP_641_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	128 
    -- CP-element group 176: 	217 
    -- CP-element group 176: 	10 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_sample_start_
      -- CP-element group 176: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Sample/$entry
      -- CP-element group 176: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Sample/crr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_568_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(176), ack => call_stmt_568_call_req_0); -- 
    initIfMaps_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(128) & initIfMaps_CP_641_elements(217) & initIfMaps_CP_641_elements(10);
      gj_initIfMaps_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_sample_completed_
      -- CP-element group 177: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Sample/$exit
      -- CP-element group 177: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Sample/cra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_568_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_568_call_ack_0, ack => initIfMaps_CP_641_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	0 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_update_completed_
      -- CP-element group 178: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Update/$exit
      -- CP-element group 178: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_568_Update/cca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:call_stmt_568_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_568_call_ack_1, ack => initIfMaps_CP_641_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	198 
    -- CP-element group 179: 	181 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	182 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_sample_start_
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/$entry
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/array_obj_ref_571_Split/$entry
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/array_obj_ref_571_Split/$exit
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/array_obj_ref_571_Split/split_req
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/array_obj_ref_571_Split/split_ack
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/$entry
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/word_0/$entry
      -- CP-element group 179: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => initIfMaps_CP_641_elements(179), ack => array_obj_ref_571_store_0_req_0); -- 
    initIfMaps_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(198) & initIfMaps_CP_641_elements(181) & initIfMaps_CP_641_elements(178);
      gj_initIfMaps_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	0 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	233 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_sample_complete
      -- CP-element group 180: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Sample/$exit
      -- CP-element group 180: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_index_offset_ack_0, ack => initIfMaps_CP_641_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	0 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (13) 
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_word_address_calculated
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_root_address_calculated
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_offset_calculated
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Update/$exit
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_final_index_sum_regn_Update/ack
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_base_plus_offset/$entry
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_base_plus_offset/$exit
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_base_plus_offset/sum_rename_req
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_base_plus_offset/sum_rename_ack
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_word_addrgen/$entry
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_word_addrgen/$exit
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_word_addrgen/root_register_req
      -- CP-element group 181: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_index_offset_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_index_offset_ack_1, ack => initIfMaps_CP_641_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_sample_completed_
      -- CP-element group 182: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/$exit
      -- CP-element group 182: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/$exit
      -- CP-element group 182: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/word_0/$exit
      -- CP-element group 182: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_store_0_ack_0, ack => initIfMaps_CP_641_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	0 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	233 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_update_completed_
      -- CP-element group 183: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/$exit
      -- CP-element group 183: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/$exit
      -- CP-element group 183: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/word_0/$exit
      -- CP-element group 183: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_571_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:array_obj_ref_571_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_store_0_ack_1, ack => initIfMaps_CP_641_elements(183)); -- 
    -- CP-element group 184:  transition  delay-element  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	35 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	43 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_304_array_obj_ref_323_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(184) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(184) is a control-delay.
    cp_element_184_delay: control_delay_element  generic map(name => " 184_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(35), ack => initIfMaps_CP_641_elements(184), clk => clk, reset =>reset);
    -- CP-element group 185:  transition  delay-element  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	44 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	52 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_323_array_obj_ref_342_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(185) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(185) is a control-delay.
    cp_element_185_delay: control_delay_element  generic map(name => " 185_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(44), ack => initIfMaps_CP_641_elements(185), clk => clk, reset =>reset);
    -- CP-element group 186:  transition  delay-element  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	53 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	61 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_342_array_obj_ref_361_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(186) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(186) is a control-delay.
    cp_element_186_delay: control_delay_element  generic map(name => " 186_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(53), ack => initIfMaps_CP_641_elements(186), clk => clk, reset =>reset);
    -- CP-element group 187:  transition  delay-element  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	62 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	70 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_361_array_obj_ref_380_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(187) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(187) is a control-delay.
    cp_element_187_delay: control_delay_element  generic map(name => " 187_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(62), ack => initIfMaps_CP_641_elements(187), clk => clk, reset =>reset);
    -- CP-element group 188:  transition  delay-element  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	71 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	79 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_380_array_obj_ref_399_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(188) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(188) is a control-delay.
    cp_element_188_delay: control_delay_element  generic map(name => " 188_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(71), ack => initIfMaps_CP_641_elements(188), clk => clk, reset =>reset);
    -- CP-element group 189:  transition  delay-element  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	80 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	88 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_399_array_obj_ref_418_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(189) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(189) is a control-delay.
    cp_element_189_delay: control_delay_element  generic map(name => " 189_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(80), ack => initIfMaps_CP_641_elements(189), clk => clk, reset =>reset);
    -- CP-element group 190:  transition  delay-element  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	89 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	97 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_418_array_obj_ref_437_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(190) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(190) is a control-delay.
    cp_element_190_delay: control_delay_element  generic map(name => " 190_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(89), ack => initIfMaps_CP_641_elements(190), clk => clk, reset =>reset);
    -- CP-element group 191:  transition  delay-element  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	98 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	106 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_437_array_obj_ref_456_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(191) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(191) is a control-delay.
    cp_element_191_delay: control_delay_element  generic map(name => " 191_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(98), ack => initIfMaps_CP_641_elements(191), clk => clk, reset =>reset);
    -- CP-element group 192:  transition  delay-element  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	107 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	112 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_456_array_obj_ref_469_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(192) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(192) is a control-delay.
    cp_element_192_delay: control_delay_element  generic map(name => " 192_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(107), ack => initIfMaps_CP_641_elements(192), clk => clk, reset =>reset);
    -- CP-element group 193:  transition  delay-element  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	113 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	118 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_469_array_obj_ref_482_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(193) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(193) is a control-delay.
    cp_element_193_delay: control_delay_element  generic map(name => " 193_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(113), ack => initIfMaps_CP_641_elements(193), clk => clk, reset =>reset);
    -- CP-element group 194:  transition  delay-element  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	119 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	124 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_482_array_obj_ref_495_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(194) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(194) is a control-delay.
    cp_element_194_delay: control_delay_element  generic map(name => " 194_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(119), ack => initIfMaps_CP_641_elements(194), clk => clk, reset =>reset);
    -- CP-element group 195:  transition  delay-element  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	125 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	145 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_495_array_obj_ref_528_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(195) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(195) is a control-delay.
    cp_element_195_delay: control_delay_element  generic map(name => " 195_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(125), ack => initIfMaps_CP_641_elements(195), clk => clk, reset =>reset);
    -- CP-element group 196:  transition  delay-element  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	148 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	158 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_528_array_obj_ref_544_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(196) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(196) is a control-delay.
    cp_element_196_delay: control_delay_element  generic map(name => " 196_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(148), ack => initIfMaps_CP_641_elements(196), clk => clk, reset =>reset);
    -- CP-element group 197:  transition  delay-element  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	161 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	171 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_544_array_obj_ref_560_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(197)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(197)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(197) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(197) is a control-delay.
    cp_element_197_delay: control_delay_element  generic map(name => " 197_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(161), ack => initIfMaps_CP_641_elements(197), clk => clk, reset =>reset);
    -- CP-element group 198:  transition  delay-element  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	174 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	179 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_560_array_obj_ref_571_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(198)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(198)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(198) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(174), ack => initIfMaps_CP_641_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  transition  delay-element  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	12 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	16 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_255_call_stmt_268_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(199)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(199)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(199) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(199) is a control-delay.
    cp_element_199_delay: control_delay_element  generic map(name => " 199_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(12), ack => initIfMaps_CP_641_elements(199), clk => clk, reset =>reset);
    -- CP-element group 200:  transition  delay-element  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	18 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	22 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_268_call_stmt_281_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(200)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(200)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(200) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(200) is a control-delay.
    cp_element_200_delay: control_delay_element  generic map(name => " 200_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(18), ack => initIfMaps_CP_641_elements(200), clk => clk, reset =>reset);
    -- CP-element group 201:  transition  delay-element  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	24 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	28 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_281_call_stmt_294_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(201)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(201)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(201) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(201) is a control-delay.
    cp_element_201_delay: control_delay_element  generic map(name => " 201_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(24), ack => initIfMaps_CP_641_elements(201), clk => clk, reset =>reset);
    -- CP-element group 202:  transition  delay-element  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	30 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	37 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_294_call_stmt_313_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(202)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(202)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(202) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(202) is a control-delay.
    cp_element_202_delay: control_delay_element  generic map(name => " 202_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(30), ack => initIfMaps_CP_641_elements(202), clk => clk, reset =>reset);
    -- CP-element group 203:  transition  delay-element  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	39 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	46 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_313_call_stmt_332_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(203)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(203)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(203) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(39), ack => initIfMaps_CP_641_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  transition  delay-element  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	48 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	55 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_332_call_stmt_351_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(204)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(204)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(204) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(204) is a control-delay.
    cp_element_204_delay: control_delay_element  generic map(name => " 204_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(48), ack => initIfMaps_CP_641_elements(204), clk => clk, reset =>reset);
    -- CP-element group 205:  transition  delay-element  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	57 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	64 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_351_call_stmt_370_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(205)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(205)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(205) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(205) is a control-delay.
    cp_element_205_delay: control_delay_element  generic map(name => " 205_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(57), ack => initIfMaps_CP_641_elements(205), clk => clk, reset =>reset);
    -- CP-element group 206:  transition  delay-element  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	66 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	73 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_370_call_stmt_389_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(206)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(206)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(206) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(206) is a control-delay.
    cp_element_206_delay: control_delay_element  generic map(name => " 206_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(66), ack => initIfMaps_CP_641_elements(206), clk => clk, reset =>reset);
    -- CP-element group 207:  transition  delay-element  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	75 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	82 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_389_call_stmt_408_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(207)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(207)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(207) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(207) is a control-delay.
    cp_element_207_delay: control_delay_element  generic map(name => " 207_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(75), ack => initIfMaps_CP_641_elements(207), clk => clk, reset =>reset);
    -- CP-element group 208:  transition  delay-element  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	84 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	91 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_408_call_stmt_427_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(208)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(208)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(208) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(208) is a control-delay.
    cp_element_208_delay: control_delay_element  generic map(name => " 208_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(84), ack => initIfMaps_CP_641_elements(208), clk => clk, reset =>reset);
    -- CP-element group 209:  transition  delay-element  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	93 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	100 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_427_call_stmt_446_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(209)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(209)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(209) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(209) is a control-delay.
    cp_element_209_delay: control_delay_element  generic map(name => " 209_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(93), ack => initIfMaps_CP_641_elements(209), clk => clk, reset =>reset);
    -- CP-element group 210:  transition  delay-element  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	102 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	109 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_446_call_stmt_465_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(210)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(210)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(210) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(210) is a control-delay.
    cp_element_210_delay: control_delay_element  generic map(name => " 210_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(102), ack => initIfMaps_CP_641_elements(210), clk => clk, reset =>reset);
    -- CP-element group 211:  transition  delay-element  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	111 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	115 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_465_call_stmt_478_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(211)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(211)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(211) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(211) is a control-delay.
    cp_element_211_delay: control_delay_element  generic map(name => " 211_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(111), ack => initIfMaps_CP_641_elements(211), clk => clk, reset =>reset);
    -- CP-element group 212:  transition  delay-element  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	117 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	121 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_478_call_stmt_491_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(212)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(212)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(212) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(212) is a control-delay.
    cp_element_212_delay: control_delay_element  generic map(name => " 212_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(117), ack => initIfMaps_CP_641_elements(212), clk => clk, reset =>reset);
    -- CP-element group 213:  transition  delay-element  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	123 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	129 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_491_call_stmt_509_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(213)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(213)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(213) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(213) is a control-delay.
    cp_element_213_delay: control_delay_element  generic map(name => " 213_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(123), ack => initIfMaps_CP_641_elements(213), clk => clk, reset =>reset);
    -- CP-element group 214:  transition  delay-element  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	131 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	137 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_509_call_stmt_520_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(214)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(214)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(214) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(214) is a control-delay.
    cp_element_214_delay: control_delay_element  generic map(name => " 214_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(131), ack => initIfMaps_CP_641_elements(214), clk => clk, reset =>reset);
    -- CP-element group 215:  transition  delay-element  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	139 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	150 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_520_call_stmt_536_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(215)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(215)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(215) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(215) is a control-delay.
    cp_element_215_delay: control_delay_element  generic map(name => " 215_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(139), ack => initIfMaps_CP_641_elements(215), clk => clk, reset =>reset);
    -- CP-element group 216:  transition  delay-element  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	152 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	163 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_536_call_stmt_552_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(216)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(216)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(216) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(216) is a control-delay.
    cp_element_216_delay: control_delay_element  generic map(name => " 216_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(152), ack => initIfMaps_CP_641_elements(216), clk => clk, reset =>reset);
    -- CP-element group 217:  transition  delay-element  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	165 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	176 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 assign_stmt_208_to_assign_stmt_577/call_stmt_552_call_stmt_568_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(217)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(217)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(217) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(217) is a control-delay.
    cp_element_217_delay: control_delay_element  generic map(name => " 217_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(165), ack => initIfMaps_CP_641_elements(217), clk => clk, reset =>reset);
    -- CP-element group 218:  transition  delay-element  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	14 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	19 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_259_array_obj_ref_272_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(218)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(218)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(218) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(218) is a control-delay.
    cp_element_218_delay: control_delay_element  generic map(name => " 218_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(14), ack => initIfMaps_CP_641_elements(218), clk => clk, reset =>reset);
    -- CP-element group 219:  transition  delay-element  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	20 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	25 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_272_array_obj_ref_285_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(219)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(219)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(219) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(219) is a control-delay.
    cp_element_219_delay: control_delay_element  generic map(name => " 219_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(20), ack => initIfMaps_CP_641_elements(219), clk => clk, reset =>reset);
    -- CP-element group 220:  transition  delay-element  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	26 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	31 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_285_array_obj_ref_298_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(220)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(220)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(220) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(220) is a control-delay.
    cp_element_220_delay: control_delay_element  generic map(name => " 220_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(26), ack => initIfMaps_CP_641_elements(220), clk => clk, reset =>reset);
    -- CP-element group 221:  transition  delay-element  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	32 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	40 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_298_array_obj_ref_317_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(221)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(221)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(221) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(221) is a control-delay.
    cp_element_221_delay: control_delay_element  generic map(name => " 221_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(32), ack => initIfMaps_CP_641_elements(221), clk => clk, reset =>reset);
    -- CP-element group 222:  transition  delay-element  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	41 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	49 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_317_array_obj_ref_336_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(222)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(222)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(222) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(222) is a control-delay.
    cp_element_222_delay: control_delay_element  generic map(name => " 222_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(41), ack => initIfMaps_CP_641_elements(222), clk => clk, reset =>reset);
    -- CP-element group 223:  transition  delay-element  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	50 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	58 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_336_array_obj_ref_355_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(223)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(223)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(223) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(223) is a control-delay.
    cp_element_223_delay: control_delay_element  generic map(name => " 223_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(50), ack => initIfMaps_CP_641_elements(223), clk => clk, reset =>reset);
    -- CP-element group 224:  transition  delay-element  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	59 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	67 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_355_array_obj_ref_374_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(224)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(224)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(224) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(224) is a control-delay.
    cp_element_224_delay: control_delay_element  generic map(name => " 224_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(59), ack => initIfMaps_CP_641_elements(224), clk => clk, reset =>reset);
    -- CP-element group 225:  transition  delay-element  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	68 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	76 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_374_array_obj_ref_393_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(225)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(225)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(225) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(225) is a control-delay.
    cp_element_225_delay: control_delay_element  generic map(name => " 225_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(68), ack => initIfMaps_CP_641_elements(225), clk => clk, reset =>reset);
    -- CP-element group 226:  transition  delay-element  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	77 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	85 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_393_array_obj_ref_412_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(226)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(226)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(226) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(226) is a control-delay.
    cp_element_226_delay: control_delay_element  generic map(name => " 226_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(77), ack => initIfMaps_CP_641_elements(226), clk => clk, reset =>reset);
    -- CP-element group 227:  transition  delay-element  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	86 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	94 
    -- CP-element group 227:  members (1) 
      -- CP-element group 227: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_412_array_obj_ref_431_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(227)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(227)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(227) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(227) is a control-delay.
    cp_element_227_delay: control_delay_element  generic map(name => " 227_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(86), ack => initIfMaps_CP_641_elements(227), clk => clk, reset =>reset);
    -- CP-element group 228:  transition  delay-element  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	95 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	103 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_431_array_obj_ref_450_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(228)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(228)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(228) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(228) is a control-delay.
    cp_element_228_delay: control_delay_element  generic map(name => " 228_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(95), ack => initIfMaps_CP_641_elements(228), clk => clk, reset =>reset);
    -- CP-element group 229:  transition  delay-element  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	104 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	132 
    -- CP-element group 229:  members (1) 
      -- CP-element group 229: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_450_array_obj_ref_512_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(229)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(229)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(229) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(229) is a control-delay.
    cp_element_229_delay: control_delay_element  generic map(name => " 229_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(104), ack => initIfMaps_CP_641_elements(229), clk => clk, reset =>reset);
    -- CP-element group 230:  transition  delay-element  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	135 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	140 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_512_array_obj_ref_523_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(230)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(230)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(230) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(230) is a control-delay.
    cp_element_230_delay: control_delay_element  generic map(name => " 230_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(135), ack => initIfMaps_CP_641_elements(230), clk => clk, reset =>reset);
    -- CP-element group 231:  transition  delay-element  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	143 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	153 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_523_array_obj_ref_539_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(231)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(231)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(231) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(231) is a control-delay.
    cp_element_231_delay: control_delay_element  generic map(name => " 231_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(143), ack => initIfMaps_CP_641_elements(231), clk => clk, reset =>reset);
    -- CP-element group 232:  transition  delay-element  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	156 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	166 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 assign_stmt_208_to_assign_stmt_577/array_obj_ref_539_array_obj_ref_555_delay
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(232)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(232)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(232) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group initIfMaps_CP_641_elements(232) is a control-delay.
    cp_element_232_delay: control_delay_element  generic map(name => " 232_delay", delay_value => 1)  port map(req => initIfMaps_CP_641_elements(156), ack => initIfMaps_CP_641_elements(232), clk => clk, reset =>reset);
    -- CP-element group 233:  join  transition  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	15 
    -- CP-element group 233: 	21 
    -- CP-element group 233: 	27 
    -- CP-element group 233: 	78 
    -- CP-element group 233: 	149 
    -- CP-element group 233: 	133 
    -- CP-element group 233: 	69 
    -- CP-element group 233: 	167 
    -- CP-element group 233: 	96 
    -- CP-element group 233: 	180 
    -- CP-element group 233: 	183 
    -- CP-element group 233: 	126 
    -- CP-element group 233: 	81 
    -- CP-element group 233: 	87 
    -- CP-element group 233: 	120 
    -- CP-element group 233: 	63 
    -- CP-element group 233: 	159 
    -- CP-element group 233: 	162 
    -- CP-element group 233: 	136 
    -- CP-element group 233: 	72 
    -- CP-element group 233: 	141 
    -- CP-element group 233: 	99 
    -- CP-element group 233: 	146 
    -- CP-element group 233: 	170 
    -- CP-element group 233: 	108 
    -- CP-element group 233: 	60 
    -- CP-element group 233: 	157 
    -- CP-element group 233: 	172 
    -- CP-element group 233: 	90 
    -- CP-element group 233: 	105 
    -- CP-element group 233: 	154 
    -- CP-element group 233: 	114 
    -- CP-element group 233: 	144 
    -- CP-element group 233: 	175 
    -- CP-element group 233: 	33 
    -- CP-element group 233: 	36 
    -- CP-element group 233: 	42 
    -- CP-element group 233: 	45 
    -- CP-element group 233: 	51 
    -- CP-element group 233: 	54 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (2) 
      -- CP-element group 233: 	 $exit
      -- CP-element group 233: 	 assign_stmt_208_to_assign_stmt_577/$exit
      -- 
    -- logger for CP element group initIfMaps_CP_641_elements(233)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and initIfMaps_CP_641_elements(233)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:initIfMaps:CP:initIfMaps_CP_641_elements(233) fired."); 
        -- 
      end if; --
    end process; 
    initIfMaps_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 39) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1);
      constant place_markings: IntegerArray(0 to 39)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0);
      constant place_delays: IntegerArray(0 to 39) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0);
      constant joinName: string(1 to 31) := "initIfMaps_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 40); -- 
    begin -- 
      preds <= initIfMaps_CP_641_elements(15) & initIfMaps_CP_641_elements(21) & initIfMaps_CP_641_elements(27) & initIfMaps_CP_641_elements(78) & initIfMaps_CP_641_elements(149) & initIfMaps_CP_641_elements(133) & initIfMaps_CP_641_elements(69) & initIfMaps_CP_641_elements(167) & initIfMaps_CP_641_elements(96) & initIfMaps_CP_641_elements(180) & initIfMaps_CP_641_elements(183) & initIfMaps_CP_641_elements(126) & initIfMaps_CP_641_elements(81) & initIfMaps_CP_641_elements(87) & initIfMaps_CP_641_elements(120) & initIfMaps_CP_641_elements(63) & initIfMaps_CP_641_elements(159) & initIfMaps_CP_641_elements(162) & initIfMaps_CP_641_elements(136) & initIfMaps_CP_641_elements(72) & initIfMaps_CP_641_elements(141) & initIfMaps_CP_641_elements(99) & initIfMaps_CP_641_elements(146) & initIfMaps_CP_641_elements(170) & initIfMaps_CP_641_elements(108) & initIfMaps_CP_641_elements(60) & initIfMaps_CP_641_elements(157) & initIfMaps_CP_641_elements(172) & initIfMaps_CP_641_elements(90) & initIfMaps_CP_641_elements(105) & initIfMaps_CP_641_elements(154) & initIfMaps_CP_641_elements(114) & initIfMaps_CP_641_elements(144) & initIfMaps_CP_641_elements(175) & initIfMaps_CP_641_elements(33) & initIfMaps_CP_641_elements(36) & initIfMaps_CP_641_elements(42) & initIfMaps_CP_641_elements(45) & initIfMaps_CP_641_elements(51) & initIfMaps_CP_641_elements(54);
      gj_initIfMaps_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 40, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => initIfMaps_CP_641_elements(233), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_501_wire : std_logic_vector(4 downto 0);
    signal ADD_u6_u6_216_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_222_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_228_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_234_wire : std_logic_vector(5 downto 0);
    signal EQ_u5_u1_202_wire : std_logic_vector(0 downto 0);
    signal J_3_503 : std_logic_vector(4 downto 0);
    signal R_col_to_be_replaced_511_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_511_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_522_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_522_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_527_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_527_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_538_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_538_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_543_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_543_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_554_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_554_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_559_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_559_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_570_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_570_scaled : std_logic_vector(3 downto 0);
    signal R_read_signal_250_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_263_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_276_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_289_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_308_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_327_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_346_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_365_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_384_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_403_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_422_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_441_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_460_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_473_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_486_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_504_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_515_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_531_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_547_wire_constant : std_logic_vector(0 downto 0);
    signal R_read_signal_563_wire_constant : std_logic_vector(0 downto 0);
    signal R_write_data_zero_253_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_266_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_279_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_292_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_311_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_330_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_349_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_368_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_387_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_406_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_425_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_444_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_463_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_476_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_489_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_507_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_518_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_534_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_550_wire_constant : std_logic_vector(15 downto 0);
    signal R_write_data_zero_566_wire_constant : std_logic_vector(15 downto 0);
    signal array_obj_ref_259_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_259_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_272_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_272_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_285_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_285_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_298_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_298_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_304_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_304_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_317_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_317_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_323_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_323_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_336_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_336_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_342_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_342_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_355_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_355_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_361_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_361_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_374_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_374_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_380_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_380_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_393_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_393_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_399_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_399_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_412_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_412_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_418_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_418_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_431_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_431_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_437_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_437_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_450_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_450_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_456_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_456_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_469_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_469_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_482_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_482_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_495_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_495_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_512_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_523_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_523_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_528_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_528_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_539_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_539_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_544_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_544_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_555_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_555_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_560_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_560_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_571_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_571_word_offset_0 : std_logic_vector(3 downto 0);
    signal checkJZero_208 : std_logic_vector(0 downto 0);
    signal col0_240 : std_logic_vector(4 downto 0);
    signal col1_244 : std_logic_vector(4 downto 0);
    signal col2_248 : std_logic_vector(4 downto 0);
    signal konst_201_wire_constant : std_logic_vector(4 downto 0);
    signal konst_215_wire_constant : std_logic_vector(5 downto 0);
    signal konst_221_wire_constant : std_logic_vector(5 downto 0);
    signal konst_227_wire_constant : std_logic_vector(5 downto 0);
    signal konst_233_wire_constant : std_logic_vector(5 downto 0);
    signal konst_500_wire_constant : std_logic_vector(4 downto 0);
    signal rdata_I00_255 : std_logic_vector(15 downto 0);
    signal rdata_I01_268 : std_logic_vector(15 downto 0);
    signal rdata_I02_281 : std_logic_vector(15 downto 0);
    signal rdata_I10_294 : std_logic_vector(15 downto 0);
    signal rdata_I11_313 : std_logic_vector(15 downto 0);
    signal rdata_I12_332 : std_logic_vector(15 downto 0);
    signal rdata_I20_351 : std_logic_vector(15 downto 0);
    signal rdata_I21_370 : std_logic_vector(15 downto 0);
    signal rdata_I22_389 : std_logic_vector(15 downto 0);
    signal rdata_I30_408 : std_logic_vector(15 downto 0);
    signal rdata_I31_427 : std_logic_vector(15 downto 0);
    signal rdata_I32_446 : std_logic_vector(15 downto 0);
    signal rdata_I40_465 : std_logic_vector(15 downto 0);
    signal rdata_I41_478 : std_logic_vector(15 downto 0);
    signal rdata_I42_491 : std_logic_vector(15 downto 0);
    signal rdata_ifmap0_509 : std_logic_vector(15 downto 0);
    signal rdata_ifmap1_520 : std_logic_vector(15 downto 0);
    signal rdata_ifmap2_536 : std_logic_vector(15 downto 0);
    signal rdata_ifmap3_552 : std_logic_vector(15 downto 0);
    signal rdata_ifmap4_568 : std_logic_vector(15 downto 0);
    signal rowI_1_218 : std_logic_vector(5 downto 0);
    signal rowI_212 : std_logic_vector(5 downto 0);
    signal rowI_2_224 : std_logic_vector(5 downto 0);
    signal rowI_3_230 : std_logic_vector(5 downto 0);
    signal rowI_4_236 : std_logic_vector(5 downto 0);
    signal type_cast_204_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_206_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_read_signal_250_wire_constant <= "1";
    R_read_signal_263_wire_constant <= "1";
    R_read_signal_276_wire_constant <= "1";
    R_read_signal_289_wire_constant <= "1";
    R_read_signal_308_wire_constant <= "1";
    R_read_signal_327_wire_constant <= "1";
    R_read_signal_346_wire_constant <= "1";
    R_read_signal_365_wire_constant <= "1";
    R_read_signal_384_wire_constant <= "1";
    R_read_signal_403_wire_constant <= "1";
    R_read_signal_422_wire_constant <= "1";
    R_read_signal_441_wire_constant <= "1";
    R_read_signal_460_wire_constant <= "1";
    R_read_signal_473_wire_constant <= "1";
    R_read_signal_486_wire_constant <= "1";
    R_read_signal_504_wire_constant <= "1";
    R_read_signal_515_wire_constant <= "1";
    R_read_signal_531_wire_constant <= "1";
    R_read_signal_547_wire_constant <= "1";
    R_read_signal_563_wire_constant <= "1";
    R_write_data_zero_253_wire_constant <= "0000000000000000";
    R_write_data_zero_266_wire_constant <= "0000000000000000";
    R_write_data_zero_279_wire_constant <= "0000000000000000";
    R_write_data_zero_292_wire_constant <= "0000000000000000";
    R_write_data_zero_311_wire_constant <= "0000000000000000";
    R_write_data_zero_330_wire_constant <= "0000000000000000";
    R_write_data_zero_349_wire_constant <= "0000000000000000";
    R_write_data_zero_368_wire_constant <= "0000000000000000";
    R_write_data_zero_387_wire_constant <= "0000000000000000";
    R_write_data_zero_406_wire_constant <= "0000000000000000";
    R_write_data_zero_425_wire_constant <= "0000000000000000";
    R_write_data_zero_444_wire_constant <= "0000000000000000";
    R_write_data_zero_463_wire_constant <= "0000000000000000";
    R_write_data_zero_476_wire_constant <= "0000000000000000";
    R_write_data_zero_489_wire_constant <= "0000000000000000";
    R_write_data_zero_507_wire_constant <= "0000000000000000";
    R_write_data_zero_518_wire_constant <= "0000000000000000";
    R_write_data_zero_534_wire_constant <= "0000000000000000";
    R_write_data_zero_550_wire_constant <= "0000000000000000";
    R_write_data_zero_566_wire_constant <= "0000000000000000";
    array_obj_ref_259_word_address_0 <= "0000";
    array_obj_ref_272_word_address_0 <= "0001";
    array_obj_ref_285_word_address_0 <= "0010";
    array_obj_ref_298_word_address_0 <= "0100";
    array_obj_ref_304_word_address_0 <= "0000";
    array_obj_ref_317_word_address_0 <= "0101";
    array_obj_ref_323_word_address_0 <= "0001";
    array_obj_ref_336_word_address_0 <= "0110";
    array_obj_ref_342_word_address_0 <= "0010";
    array_obj_ref_355_word_address_0 <= "1000";
    array_obj_ref_361_word_address_0 <= "0100";
    array_obj_ref_374_word_address_0 <= "1001";
    array_obj_ref_380_word_address_0 <= "0101";
    array_obj_ref_393_word_address_0 <= "1010";
    array_obj_ref_399_word_address_0 <= "0110";
    array_obj_ref_412_word_address_0 <= "1100";
    array_obj_ref_418_word_address_0 <= "1000";
    array_obj_ref_431_word_address_0 <= "1101";
    array_obj_ref_437_word_address_0 <= "1001";
    array_obj_ref_450_word_address_0 <= "1110";
    array_obj_ref_456_word_address_0 <= "1010";
    array_obj_ref_469_word_address_0 <= "1100";
    array_obj_ref_482_word_address_0 <= "1101";
    array_obj_ref_495_word_address_0 <= "1110";
    array_obj_ref_512_constant_part_of_offset <= "0000";
    array_obj_ref_512_offset_scale_factor_0 <= "0100";
    array_obj_ref_512_offset_scale_factor_1 <= "0001";
    array_obj_ref_512_resized_base_address <= "0000";
    array_obj_ref_512_word_offset_0 <= "0000";
    array_obj_ref_523_constant_part_of_offset <= "0100";
    array_obj_ref_523_offset_scale_factor_0 <= "0100";
    array_obj_ref_523_offset_scale_factor_1 <= "0001";
    array_obj_ref_523_resized_base_address <= "0000";
    array_obj_ref_523_word_offset_0 <= "0000";
    array_obj_ref_528_constant_part_of_offset <= "0000";
    array_obj_ref_528_offset_scale_factor_0 <= "0100";
    array_obj_ref_528_offset_scale_factor_1 <= "0001";
    array_obj_ref_528_resized_base_address <= "0000";
    array_obj_ref_528_word_offset_0 <= "0000";
    array_obj_ref_539_constant_part_of_offset <= "1000";
    array_obj_ref_539_offset_scale_factor_0 <= "0100";
    array_obj_ref_539_offset_scale_factor_1 <= "0001";
    array_obj_ref_539_resized_base_address <= "0000";
    array_obj_ref_539_word_offset_0 <= "0000";
    array_obj_ref_544_constant_part_of_offset <= "0100";
    array_obj_ref_544_offset_scale_factor_0 <= "0100";
    array_obj_ref_544_offset_scale_factor_1 <= "0001";
    array_obj_ref_544_resized_base_address <= "0000";
    array_obj_ref_544_word_offset_0 <= "0000";
    array_obj_ref_555_constant_part_of_offset <= "1100";
    array_obj_ref_555_offset_scale_factor_0 <= "0100";
    array_obj_ref_555_offset_scale_factor_1 <= "0001";
    array_obj_ref_555_resized_base_address <= "0000";
    array_obj_ref_555_word_offset_0 <= "0000";
    array_obj_ref_560_constant_part_of_offset <= "1000";
    array_obj_ref_560_offset_scale_factor_0 <= "0100";
    array_obj_ref_560_offset_scale_factor_1 <= "0001";
    array_obj_ref_560_resized_base_address <= "0000";
    array_obj_ref_560_word_offset_0 <= "0000";
    array_obj_ref_571_constant_part_of_offset <= "1100";
    array_obj_ref_571_offset_scale_factor_0 <= "0100";
    array_obj_ref_571_offset_scale_factor_1 <= "0001";
    array_obj_ref_571_resized_base_address <= "0000";
    array_obj_ref_571_word_offset_0 <= "0000";
    col0_240 <= "00000";
    col1_244 <= "00001";
    col2_248 <= "00010";
    konst_201_wire_constant <= "00000";
    konst_215_wire_constant <= "000001";
    konst_221_wire_constant <= "000010";
    konst_227_wire_constant <= "000011";
    konst_233_wire_constant <= "000100";
    konst_500_wire_constant <= "00011";
    type_cast_204_wire_constant <= "0";
    type_cast_206_wire_constant <= "1";
    -- logger for split-operator MUX_207_inst flow-through 
    process(checkJZero_208) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:MUX_207_inst:flowthrough inputs: " & " EQ_u5_u1_202_wire = "& Convert_SLV_To_Hex_String(EQ_u5_u1_202_wire) & " type_cast_204_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_204_wire_constant) & " type_cast_206_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_206_wire_constant) & " outputs:" & " checkJZero_208= "  & Convert_SLV_To_Hex_String(checkJZero_208));
      --
    end process; 
    -- flow-through select operator MUX_207_inst
    checkJZero_208 <= type_cast_204_wire_constant when (EQ_u5_u1_202_wire(0) /=  '0') else type_cast_206_wire_constant;
    -- logger for split-operator type_cast_211_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_211_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_211_inst:started:   inputs: " & " I_buffer = "& Convert_SLV_To_Hex_String(I_buffer));
          --
        end if; 
        if type_cast_211_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_211_inst:finished:  outputs: " & " rowI_212= "  & Convert_SLV_To_Hex_String(rowI_212));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_211_inst_req_0;
      type_cast_211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_211_inst_req_1;
      type_cast_211_inst_ack_1<= rack(0);
      type_cast_211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => I_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowI_212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_217_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_217_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_217_inst:started:   inputs: " & " ADD_u6_u6_216_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_216_wire));
          --
        end if; 
        if type_cast_217_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_217_inst:finished:  outputs: " & " rowI_1_218= "  & Convert_SLV_To_Hex_String(rowI_1_218));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_217_inst_req_0;
      type_cast_217_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_217_inst_req_1;
      type_cast_217_inst_ack_1<= rack(0);
      type_cast_217_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_217_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u6_u6_216_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowI_1_218,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_223_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_223_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_223_inst:started:   inputs: " & " ADD_u6_u6_222_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_222_wire));
          --
        end if; 
        if type_cast_223_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_223_inst:finished:  outputs: " & " rowI_2_224= "  & Convert_SLV_To_Hex_String(rowI_2_224));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_223_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_223_inst_req_0;
      type_cast_223_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_223_inst_req_1;
      type_cast_223_inst_ack_1<= rack(0);
      type_cast_223_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_223_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u6_u6_222_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowI_2_224,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_229_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_229_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_229_inst:started:   inputs: " & " ADD_u6_u6_228_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_228_wire));
          --
        end if; 
        if type_cast_229_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_229_inst:finished:  outputs: " & " rowI_3_230= "  & Convert_SLV_To_Hex_String(rowI_3_230));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_229_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_229_inst_req_0;
      type_cast_229_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_229_inst_req_1;
      type_cast_229_inst_ack_1<= rack(0);
      type_cast_229_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_229_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u6_u6_228_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowI_3_230,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_235_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_235_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_235_inst:started:   inputs: " & " ADD_u6_u6_234_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_234_wire));
          --
        end if; 
        if type_cast_235_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_235_inst:finished:  outputs: " & " rowI_4_236= "  & Convert_SLV_To_Hex_String(rowI_4_236));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_235_inst_req_0;
      type_cast_235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_235_inst_req_1;
      type_cast_235_inst_ack_1<= rack(0);
      type_cast_235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u6_u6_234_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowI_4_236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_502_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_502_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_502_inst:started:   inputs: " & " ADD_u5_u5_501_wire = "& Convert_SLV_To_Hex_String(ADD_u5_u5_501_wire));
          --
        end if; 
        if type_cast_502_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:type_cast_502_inst:finished:  outputs: " & " J_3_503= "  & Convert_SLV_To_Hex_String(J_3_503));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_502_inst_req_0;
      type_cast_502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_502_inst_req_1;
      type_cast_502_inst_ack_1<= rack(0);
      type_cast_502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 5,
        out_data_width => 5,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u5_u5_501_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => J_3_503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_259_gather_scatter flow-through 
    process(array_obj_ref_259_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_259_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I00_255 = "& Convert_SLV_To_Hex_String(rdata_I00_255) & "outputs: " & " array_obj_ref_259_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_259_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_259_gather_scatter
    process(rdata_I00_255) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I00_255;
      ov(15 downto 0) := iv;
      array_obj_ref_259_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_272_gather_scatter flow-through 
    process(array_obj_ref_272_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_272_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I01_268 = "& Convert_SLV_To_Hex_String(rdata_I01_268) & "outputs: " & " array_obj_ref_272_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_272_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_272_gather_scatter
    process(rdata_I01_268) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I01_268;
      ov(15 downto 0) := iv;
      array_obj_ref_272_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_285_gather_scatter flow-through 
    process(array_obj_ref_285_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_285_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I02_281 = "& Convert_SLV_To_Hex_String(rdata_I02_281) & "outputs: " & " array_obj_ref_285_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_285_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_285_gather_scatter
    process(rdata_I02_281) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I02_281;
      ov(15 downto 0) := iv;
      array_obj_ref_285_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_298_gather_scatter flow-through 
    process(array_obj_ref_298_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_298_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I10_294 = "& Convert_SLV_To_Hex_String(rdata_I10_294) & "outputs: " & " array_obj_ref_298_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_298_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_298_gather_scatter
    process(rdata_I10_294) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I10_294;
      ov(15 downto 0) := iv;
      array_obj_ref_298_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_304_gather_scatter flow-through 
    process(array_obj_ref_304_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_304_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I10_294 = "& Convert_SLV_To_Hex_String(rdata_I10_294) & "outputs: " & " array_obj_ref_304_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_304_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_304_gather_scatter
    process(rdata_I10_294) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I10_294;
      ov(15 downto 0) := iv;
      array_obj_ref_304_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_317_gather_scatter flow-through 
    process(array_obj_ref_317_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_317_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I11_313 = "& Convert_SLV_To_Hex_String(rdata_I11_313) & "outputs: " & " array_obj_ref_317_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_317_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_317_gather_scatter
    process(rdata_I11_313) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I11_313;
      ov(15 downto 0) := iv;
      array_obj_ref_317_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_323_gather_scatter flow-through 
    process(array_obj_ref_323_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_323_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I11_313 = "& Convert_SLV_To_Hex_String(rdata_I11_313) & "outputs: " & " array_obj_ref_323_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_323_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_323_gather_scatter
    process(rdata_I11_313) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I11_313;
      ov(15 downto 0) := iv;
      array_obj_ref_323_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_336_gather_scatter flow-through 
    process(array_obj_ref_336_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_336_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I12_332 = "& Convert_SLV_To_Hex_String(rdata_I12_332) & "outputs: " & " array_obj_ref_336_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_336_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_336_gather_scatter
    process(rdata_I12_332) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I12_332;
      ov(15 downto 0) := iv;
      array_obj_ref_336_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_342_gather_scatter flow-through 
    process(array_obj_ref_342_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_342_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I12_332 = "& Convert_SLV_To_Hex_String(rdata_I12_332) & "outputs: " & " array_obj_ref_342_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_342_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_342_gather_scatter
    process(rdata_I12_332) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I12_332;
      ov(15 downto 0) := iv;
      array_obj_ref_342_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_355_gather_scatter flow-through 
    process(array_obj_ref_355_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_355_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I20_351 = "& Convert_SLV_To_Hex_String(rdata_I20_351) & "outputs: " & " array_obj_ref_355_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_355_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_355_gather_scatter
    process(rdata_I20_351) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I20_351;
      ov(15 downto 0) := iv;
      array_obj_ref_355_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_361_gather_scatter flow-through 
    process(array_obj_ref_361_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_361_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I20_351 = "& Convert_SLV_To_Hex_String(rdata_I20_351) & "outputs: " & " array_obj_ref_361_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_361_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_361_gather_scatter
    process(rdata_I20_351) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I20_351;
      ov(15 downto 0) := iv;
      array_obj_ref_361_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_374_gather_scatter flow-through 
    process(array_obj_ref_374_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_374_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I21_370 = "& Convert_SLV_To_Hex_String(rdata_I21_370) & "outputs: " & " array_obj_ref_374_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_374_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_374_gather_scatter
    process(rdata_I21_370) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I21_370;
      ov(15 downto 0) := iv;
      array_obj_ref_374_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_380_gather_scatter flow-through 
    process(array_obj_ref_380_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_380_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I21_370 = "& Convert_SLV_To_Hex_String(rdata_I21_370) & "outputs: " & " array_obj_ref_380_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_380_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_380_gather_scatter
    process(rdata_I21_370) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I21_370;
      ov(15 downto 0) := iv;
      array_obj_ref_380_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_393_gather_scatter flow-through 
    process(array_obj_ref_393_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_393_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I22_389 = "& Convert_SLV_To_Hex_String(rdata_I22_389) & "outputs: " & " array_obj_ref_393_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_393_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_393_gather_scatter
    process(rdata_I22_389) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I22_389;
      ov(15 downto 0) := iv;
      array_obj_ref_393_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_399_gather_scatter flow-through 
    process(array_obj_ref_399_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_399_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I22_389 = "& Convert_SLV_To_Hex_String(rdata_I22_389) & "outputs: " & " array_obj_ref_399_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_399_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_399_gather_scatter
    process(rdata_I22_389) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I22_389;
      ov(15 downto 0) := iv;
      array_obj_ref_399_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_412_gather_scatter flow-through 
    process(array_obj_ref_412_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_412_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I30_408 = "& Convert_SLV_To_Hex_String(rdata_I30_408) & "outputs: " & " array_obj_ref_412_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_412_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_412_gather_scatter
    process(rdata_I30_408) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I30_408;
      ov(15 downto 0) := iv;
      array_obj_ref_412_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_418_gather_scatter flow-through 
    process(array_obj_ref_418_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_418_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I30_408 = "& Convert_SLV_To_Hex_String(rdata_I30_408) & "outputs: " & " array_obj_ref_418_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_418_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_418_gather_scatter
    process(rdata_I30_408) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I30_408;
      ov(15 downto 0) := iv;
      array_obj_ref_418_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_431_gather_scatter flow-through 
    process(array_obj_ref_431_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_431_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I31_427 = "& Convert_SLV_To_Hex_String(rdata_I31_427) & "outputs: " & " array_obj_ref_431_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_431_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_431_gather_scatter
    process(rdata_I31_427) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I31_427;
      ov(15 downto 0) := iv;
      array_obj_ref_431_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_437_gather_scatter flow-through 
    process(array_obj_ref_437_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_437_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I31_427 = "& Convert_SLV_To_Hex_String(rdata_I31_427) & "outputs: " & " array_obj_ref_437_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_437_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_437_gather_scatter
    process(rdata_I31_427) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I31_427;
      ov(15 downto 0) := iv;
      array_obj_ref_437_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_450_gather_scatter flow-through 
    process(array_obj_ref_450_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_450_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I32_446 = "& Convert_SLV_To_Hex_String(rdata_I32_446) & "outputs: " & " array_obj_ref_450_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_450_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_450_gather_scatter
    process(rdata_I32_446) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I32_446;
      ov(15 downto 0) := iv;
      array_obj_ref_450_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_456_gather_scatter flow-through 
    process(array_obj_ref_456_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_456_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I32_446 = "& Convert_SLV_To_Hex_String(rdata_I32_446) & "outputs: " & " array_obj_ref_456_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_456_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_456_gather_scatter
    process(rdata_I32_446) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I32_446;
      ov(15 downto 0) := iv;
      array_obj_ref_456_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_469_gather_scatter flow-through 
    process(array_obj_ref_469_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_469_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I40_465 = "& Convert_SLV_To_Hex_String(rdata_I40_465) & "outputs: " & " array_obj_ref_469_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_469_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_469_gather_scatter
    process(rdata_I40_465) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I40_465;
      ov(15 downto 0) := iv;
      array_obj_ref_469_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_482_gather_scatter flow-through 
    process(array_obj_ref_482_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_482_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I41_478 = "& Convert_SLV_To_Hex_String(rdata_I41_478) & "outputs: " & " array_obj_ref_482_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_482_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_482_gather_scatter
    process(rdata_I41_478) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I41_478;
      ov(15 downto 0) := iv;
      array_obj_ref_482_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_495_gather_scatter flow-through 
    process(array_obj_ref_495_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_495_gather_scatter:flowthrough  inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " rdata_I42_491 = "& Convert_SLV_To_Hex_String(rdata_I42_491) & "outputs: " & " array_obj_ref_495_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_495_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_495_gather_scatter
    process(rdata_I42_491) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_I42_491;
      ov(15 downto 0) := iv;
      array_obj_ref_495_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_512_addr_0 flow-through 
    process(array_obj_ref_512_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_addr_0:flowthrough  inputs: " & " array_obj_ref_512_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_512_root_address) & "outputs: " & " array_obj_ref_512_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_512_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_512_addr_0
    process(array_obj_ref_512_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_512_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_512_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_512_gather_scatter flow-through 
    process(array_obj_ref_512_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_gather_scatter:flowthrough  inputs: " & " rdata_ifmap0_509 = "& Convert_SLV_To_Hex_String(rdata_ifmap0_509) & "outputs: " & " array_obj_ref_512_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_512_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_512_gather_scatter
    process(rdata_ifmap0_509) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap0_509;
      ov(15 downto 0) := iv;
      array_obj_ref_512_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_512_index_1_rename flow-through 
    process(R_col_to_be_replaced_511_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_511_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_511_resized) & "outputs: " & " R_col_to_be_replaced_511_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_511_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_512_index_1_rename
    process(R_col_to_be_replaced_511_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_511_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_511_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_512_index_1_resize flow-through 
    process(R_col_to_be_replaced_511_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_511_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_511_resized));
      --
    end process; 
    -- equivalence array_obj_ref_512_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_511_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_512_root_address_inst flow-through 
    process(array_obj_ref_512_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_root_address_inst:flowthrough  inputs: " & " array_obj_ref_512_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_512_final_offset) & "outputs: " & " array_obj_ref_512_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_512_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_512_root_address_inst
    process(array_obj_ref_512_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_512_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_512_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_523_addr_0 flow-through 
    process(array_obj_ref_523_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_addr_0:flowthrough  inputs: " & " array_obj_ref_523_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_523_root_address) & "outputs: " & " array_obj_ref_523_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_523_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_523_addr_0
    process(array_obj_ref_523_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_523_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_523_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_523_gather_scatter flow-through 
    process(array_obj_ref_523_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_gather_scatter:flowthrough  inputs: " & " rdata_ifmap1_520 = "& Convert_SLV_To_Hex_String(rdata_ifmap1_520) & "outputs: " & " array_obj_ref_523_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_523_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_523_gather_scatter
    process(rdata_ifmap1_520) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap1_520;
      ov(15 downto 0) := iv;
      array_obj_ref_523_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_523_index_1_rename flow-through 
    process(R_col_to_be_replaced_522_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_522_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_522_resized) & "outputs: " & " R_col_to_be_replaced_522_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_522_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_523_index_1_rename
    process(R_col_to_be_replaced_522_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_522_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_522_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_523_index_1_resize flow-through 
    process(R_col_to_be_replaced_522_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_522_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_522_resized));
      --
    end process; 
    -- equivalence array_obj_ref_523_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_522_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_523_root_address_inst flow-through 
    process(array_obj_ref_523_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_root_address_inst:flowthrough  inputs: " & " array_obj_ref_523_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_523_final_offset) & "outputs: " & " array_obj_ref_523_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_523_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_523_root_address_inst
    process(array_obj_ref_523_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_523_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_523_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_528_addr_0 flow-through 
    process(array_obj_ref_528_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_addr_0:flowthrough  inputs: " & " array_obj_ref_528_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_528_root_address) & "outputs: " & " array_obj_ref_528_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_528_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_528_addr_0
    process(array_obj_ref_528_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_528_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_528_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_528_gather_scatter flow-through 
    process(array_obj_ref_528_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_gather_scatter:flowthrough  inputs: " & " rdata_ifmap1_520 = "& Convert_SLV_To_Hex_String(rdata_ifmap1_520) & "outputs: " & " array_obj_ref_528_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_528_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_528_gather_scatter
    process(rdata_ifmap1_520) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap1_520;
      ov(15 downto 0) := iv;
      array_obj_ref_528_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_528_index_1_rename flow-through 
    process(R_col_to_be_replaced_527_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_527_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_527_resized) & "outputs: " & " R_col_to_be_replaced_527_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_527_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_528_index_1_rename
    process(R_col_to_be_replaced_527_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_527_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_527_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_528_index_1_resize flow-through 
    process(R_col_to_be_replaced_527_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_527_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_527_resized));
      --
    end process; 
    -- equivalence array_obj_ref_528_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_527_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_528_root_address_inst flow-through 
    process(array_obj_ref_528_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_root_address_inst:flowthrough  inputs: " & " array_obj_ref_528_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_528_final_offset) & "outputs: " & " array_obj_ref_528_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_528_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_528_root_address_inst
    process(array_obj_ref_528_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_528_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_528_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_539_addr_0 flow-through 
    process(array_obj_ref_539_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_addr_0:flowthrough  inputs: " & " array_obj_ref_539_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_539_root_address) & "outputs: " & " array_obj_ref_539_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_539_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_539_addr_0
    process(array_obj_ref_539_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_539_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_539_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_539_gather_scatter flow-through 
    process(array_obj_ref_539_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_gather_scatter:flowthrough  inputs: " & " rdata_ifmap2_536 = "& Convert_SLV_To_Hex_String(rdata_ifmap2_536) & "outputs: " & " array_obj_ref_539_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_539_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_539_gather_scatter
    process(rdata_ifmap2_536) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap2_536;
      ov(15 downto 0) := iv;
      array_obj_ref_539_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_539_index_1_rename flow-through 
    process(R_col_to_be_replaced_538_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_538_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_538_resized) & "outputs: " & " R_col_to_be_replaced_538_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_538_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_539_index_1_rename
    process(R_col_to_be_replaced_538_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_538_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_538_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_539_index_1_resize flow-through 
    process(R_col_to_be_replaced_538_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_538_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_538_resized));
      --
    end process; 
    -- equivalence array_obj_ref_539_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_538_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_539_root_address_inst flow-through 
    process(array_obj_ref_539_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_root_address_inst:flowthrough  inputs: " & " array_obj_ref_539_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_539_final_offset) & "outputs: " & " array_obj_ref_539_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_539_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_539_root_address_inst
    process(array_obj_ref_539_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_539_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_539_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_544_addr_0 flow-through 
    process(array_obj_ref_544_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_addr_0:flowthrough  inputs: " & " array_obj_ref_544_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_544_root_address) & "outputs: " & " array_obj_ref_544_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_544_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_544_addr_0
    process(array_obj_ref_544_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_544_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_544_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_544_gather_scatter flow-through 
    process(array_obj_ref_544_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_gather_scatter:flowthrough  inputs: " & " rdata_ifmap2_536 = "& Convert_SLV_To_Hex_String(rdata_ifmap2_536) & "outputs: " & " array_obj_ref_544_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_544_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_544_gather_scatter
    process(rdata_ifmap2_536) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap2_536;
      ov(15 downto 0) := iv;
      array_obj_ref_544_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_544_index_1_rename flow-through 
    process(R_col_to_be_replaced_543_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_543_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_543_resized) & "outputs: " & " R_col_to_be_replaced_543_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_543_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_544_index_1_rename
    process(R_col_to_be_replaced_543_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_543_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_543_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_544_index_1_resize flow-through 
    process(R_col_to_be_replaced_543_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_543_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_543_resized));
      --
    end process; 
    -- equivalence array_obj_ref_544_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_543_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_544_root_address_inst flow-through 
    process(array_obj_ref_544_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_root_address_inst:flowthrough  inputs: " & " array_obj_ref_544_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_544_final_offset) & "outputs: " & " array_obj_ref_544_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_544_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_544_root_address_inst
    process(array_obj_ref_544_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_544_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_544_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_555_addr_0 flow-through 
    process(array_obj_ref_555_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_addr_0:flowthrough  inputs: " & " array_obj_ref_555_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_555_root_address) & "outputs: " & " array_obj_ref_555_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_555_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_555_addr_0
    process(array_obj_ref_555_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_555_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_555_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_555_gather_scatter flow-through 
    process(array_obj_ref_555_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_gather_scatter:flowthrough  inputs: " & " rdata_ifmap3_552 = "& Convert_SLV_To_Hex_String(rdata_ifmap3_552) & "outputs: " & " array_obj_ref_555_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_555_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_555_gather_scatter
    process(rdata_ifmap3_552) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap3_552;
      ov(15 downto 0) := iv;
      array_obj_ref_555_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_555_index_1_rename flow-through 
    process(R_col_to_be_replaced_554_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_554_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_554_resized) & "outputs: " & " R_col_to_be_replaced_554_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_554_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_555_index_1_rename
    process(R_col_to_be_replaced_554_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_554_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_554_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_555_index_1_resize flow-through 
    process(R_col_to_be_replaced_554_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_554_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_554_resized));
      --
    end process; 
    -- equivalence array_obj_ref_555_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_554_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_555_root_address_inst flow-through 
    process(array_obj_ref_555_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_root_address_inst:flowthrough  inputs: " & " array_obj_ref_555_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_555_final_offset) & "outputs: " & " array_obj_ref_555_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_555_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_555_root_address_inst
    process(array_obj_ref_555_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_555_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_555_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_560_addr_0 flow-through 
    process(array_obj_ref_560_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_addr_0:flowthrough  inputs: " & " array_obj_ref_560_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_560_root_address) & "outputs: " & " array_obj_ref_560_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_560_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_560_addr_0
    process(array_obj_ref_560_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_560_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_560_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_560_gather_scatter flow-through 
    process(array_obj_ref_560_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_gather_scatter:flowthrough  inputs: " & " rdata_ifmap3_552 = "& Convert_SLV_To_Hex_String(rdata_ifmap3_552) & "outputs: " & " array_obj_ref_560_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_560_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_560_gather_scatter
    process(rdata_ifmap3_552) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap3_552;
      ov(15 downto 0) := iv;
      array_obj_ref_560_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_560_index_1_rename flow-through 
    process(R_col_to_be_replaced_559_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_559_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_559_resized) & "outputs: " & " R_col_to_be_replaced_559_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_559_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_560_index_1_rename
    process(R_col_to_be_replaced_559_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_559_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_559_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_560_index_1_resize flow-through 
    process(R_col_to_be_replaced_559_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_559_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_559_resized));
      --
    end process; 
    -- equivalence array_obj_ref_560_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_559_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_560_root_address_inst flow-through 
    process(array_obj_ref_560_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_root_address_inst:flowthrough  inputs: " & " array_obj_ref_560_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_560_final_offset) & "outputs: " & " array_obj_ref_560_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_560_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_560_root_address_inst
    process(array_obj_ref_560_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_560_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_560_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_571_addr_0 flow-through 
    process(array_obj_ref_571_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_addr_0:flowthrough  inputs: " & " array_obj_ref_571_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_571_root_address) & "outputs: " & " array_obj_ref_571_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_571_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_571_addr_0
    process(array_obj_ref_571_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_571_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_571_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_571_gather_scatter flow-through 
    process(array_obj_ref_571_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_gather_scatter:flowthrough  inputs: " & " rdata_ifmap4_568 = "& Convert_SLV_To_Hex_String(rdata_ifmap4_568) & "outputs: " & " array_obj_ref_571_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_571_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_571_gather_scatter
    process(rdata_ifmap4_568) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := rdata_ifmap4_568;
      ov(15 downto 0) := iv;
      array_obj_ref_571_data_0 <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_571_index_1_rename flow-through 
    process(R_col_to_be_replaced_570_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_570_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_570_resized) & "outputs: " & " R_col_to_be_replaced_570_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_570_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_571_index_1_rename
    process(R_col_to_be_replaced_570_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_570_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_570_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_571_index_1_resize flow-through 
    process(R_col_to_be_replaced_570_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_570_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_570_resized));
      --
    end process; 
    -- equivalence array_obj_ref_571_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_570_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_571_root_address_inst flow-through 
    process(array_obj_ref_571_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_root_address_inst:flowthrough  inputs: " & " array_obj_ref_571_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_571_final_offset) & "outputs: " & " array_obj_ref_571_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_571_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_571_root_address_inst
    process(array_obj_ref_571_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_571_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_571_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u5_u5_501_inst flow-through 
    process(ADD_u5_u5_501_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:ADD_u5_u5_501_inst:flowthrough inputs: " & " J_buffer = "& Convert_SLV_To_Hex_String(J_buffer) & " konst_500_wire_constant = "& Convert_SLV_To_Hex_String(konst_500_wire_constant) & " outputs:" & " ADD_u5_u5_501_wire= "  & Convert_SLV_To_Hex_String(ADD_u5_u5_501_wire));
      --
    end process; 
    -- binary operator ADD_u5_u5_501_inst
    process(J_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntAdd_proc(J_buffer, konst_500_wire_constant, tmp_var);
      ADD_u5_u5_501_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_216_inst flow-through 
    process(ADD_u6_u6_216_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:ADD_u6_u6_216_inst:flowthrough inputs: " & " I_buffer = "& Convert_SLV_To_Hex_String(I_buffer) & " konst_215_wire_constant = "& Convert_SLV_To_Hex_String(konst_215_wire_constant) & " outputs:" & " ADD_u6_u6_216_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_216_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_216_inst
    process(I_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_buffer, konst_215_wire_constant, tmp_var);
      ADD_u6_u6_216_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_222_inst flow-through 
    process(ADD_u6_u6_222_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:ADD_u6_u6_222_inst:flowthrough inputs: " & " I_buffer = "& Convert_SLV_To_Hex_String(I_buffer) & " konst_221_wire_constant = "& Convert_SLV_To_Hex_String(konst_221_wire_constant) & " outputs:" & " ADD_u6_u6_222_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_222_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_222_inst
    process(I_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_buffer, konst_221_wire_constant, tmp_var);
      ADD_u6_u6_222_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_228_inst flow-through 
    process(ADD_u6_u6_228_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:ADD_u6_u6_228_inst:flowthrough inputs: " & " I_buffer = "& Convert_SLV_To_Hex_String(I_buffer) & " konst_227_wire_constant = "& Convert_SLV_To_Hex_String(konst_227_wire_constant) & " outputs:" & " ADD_u6_u6_228_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_228_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_228_inst
    process(I_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_buffer, konst_227_wire_constant, tmp_var);
      ADD_u6_u6_228_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_234_inst flow-through 
    process(ADD_u6_u6_234_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:ADD_u6_u6_234_inst:flowthrough inputs: " & " I_buffer = "& Convert_SLV_To_Hex_String(I_buffer) & " konst_233_wire_constant = "& Convert_SLV_To_Hex_String(konst_233_wire_constant) & " outputs:" & " ADD_u6_u6_234_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_234_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_234_inst
    process(I_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_buffer, konst_233_wire_constant, tmp_var);
      ADD_u6_u6_234_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u5_u1_202_inst flow-through 
    process(EQ_u5_u1_202_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:EQ_u5_u1_202_inst:flowthrough inputs: " & " J_buffer = "& Convert_SLV_To_Hex_String(J_buffer) & " konst_201_wire_constant = "& Convert_SLV_To_Hex_String(konst_201_wire_constant) & " outputs:" & " EQ_u5_u1_202_wire= "  & Convert_SLV_To_Hex_String(EQ_u5_u1_202_wire));
      --
    end process; 
    -- binary operator EQ_u5_u1_202_inst
    process(J_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(J_buffer, konst_201_wire_constant, tmp_var);
      EQ_u5_u1_202_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_512_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_512_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_index_offset:started:   inputs: " & " R_col_to_be_replaced_511_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_511_scaled) & " array_obj_ref_512_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_512_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_512_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_index_offset:finished:  outputs: " & " array_obj_ref_512_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_512_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (6) : array_obj_ref_512_index_offset 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_511_scaled;
      array_obj_ref_512_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_512_index_offset_req_0;
      array_obj_ref_512_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_512_index_offset_req_1;
      array_obj_ref_512_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- logger for split-operator array_obj_ref_523_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_523_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_index_offset:started:   inputs: " & " R_col_to_be_replaced_522_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_522_scaled) & " array_obj_ref_523_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_523_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_523_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_index_offset:finished:  outputs: " & " array_obj_ref_523_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_523_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (7) : array_obj_ref_523_index_offset 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_522_scaled;
      array_obj_ref_523_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_523_index_offset_req_0;
      array_obj_ref_523_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_523_index_offset_req_1;
      array_obj_ref_523_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_7_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- logger for split-operator array_obj_ref_528_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_528_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_index_offset:started:   inputs: " & " R_col_to_be_replaced_527_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_527_scaled) & " array_obj_ref_528_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_528_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_528_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_index_offset:finished:  outputs: " & " array_obj_ref_528_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_528_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (8) : array_obj_ref_528_index_offset 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_527_scaled;
      array_obj_ref_528_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_528_index_offset_req_0;
      array_obj_ref_528_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_528_index_offset_req_1;
      array_obj_ref_528_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_8_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- logger for split-operator array_obj_ref_539_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_539_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_index_offset:started:   inputs: " & " R_col_to_be_replaced_538_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_538_scaled) & " array_obj_ref_539_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_539_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_539_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_index_offset:finished:  outputs: " & " array_obj_ref_539_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_539_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (9) : array_obj_ref_539_index_offset 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_538_scaled;
      array_obj_ref_539_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_539_index_offset_req_0;
      array_obj_ref_539_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_539_index_offset_req_1;
      array_obj_ref_539_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_9_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- logger for split-operator array_obj_ref_544_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_544_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_index_offset:started:   inputs: " & " R_col_to_be_replaced_543_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_543_scaled) & " array_obj_ref_544_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_544_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_544_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_index_offset:finished:  outputs: " & " array_obj_ref_544_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_544_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (10) : array_obj_ref_544_index_offset 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_543_scaled;
      array_obj_ref_544_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_544_index_offset_req_0;
      array_obj_ref_544_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_544_index_offset_req_1;
      array_obj_ref_544_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_10_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- logger for split-operator array_obj_ref_555_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_555_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_index_offset:started:   inputs: " & " R_col_to_be_replaced_554_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_554_scaled) & " array_obj_ref_555_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_555_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_555_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_index_offset:finished:  outputs: " & " array_obj_ref_555_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_555_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (11) : array_obj_ref_555_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_554_scaled;
      array_obj_ref_555_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_555_index_offset_req_0;
      array_obj_ref_555_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_555_index_offset_req_1;
      array_obj_ref_555_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- logger for split-operator array_obj_ref_560_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_560_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_index_offset:started:   inputs: " & " R_col_to_be_replaced_559_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_559_scaled) & " array_obj_ref_560_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_560_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_560_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_index_offset:finished:  outputs: " & " array_obj_ref_560_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_560_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (12) : array_obj_ref_560_index_offset 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_559_scaled;
      array_obj_ref_560_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_560_index_offset_req_0;
      array_obj_ref_560_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_560_index_offset_req_1;
      array_obj_ref_560_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_12_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- logger for split-operator array_obj_ref_571_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_571_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_index_offset:started:   inputs: " & " R_col_to_be_replaced_570_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_570_scaled) & " array_obj_ref_571_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_571_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_571_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_index_offset:finished:  outputs: " & " array_obj_ref_571_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_571_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (13) : array_obj_ref_571_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_570_scaled;
      array_obj_ref_571_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_571_index_offset_req_0;
      array_obj_ref_571_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_571_index_offset_req_1;
      array_obj_ref_571_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- logger for split-operator array_obj_ref_285_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_285_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_285_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_285_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_285_word_address_0) & " array_obj_ref_285_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_285_data_0));
          --
        end if; 
        if array_obj_ref_285_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_285_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_539_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_539_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_store_0:started:   inputs: " & " array_obj_ref_539_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_539_word_address_0) & " array_obj_ref_539_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_539_data_0));
          --
        end if; 
        if array_obj_ref_539_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_539_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_272_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_272_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_272_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_272_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_272_word_address_0) & " array_obj_ref_272_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_272_data_0));
          --
        end if; 
        if array_obj_ref_272_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_272_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_523_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_523_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_store_0:started:   inputs: " & " array_obj_ref_523_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_523_word_address_0) & " array_obj_ref_523_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_523_data_0));
          --
        end if; 
        if array_obj_ref_523_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_523_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_259_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_259_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_259_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_259_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_259_word_address_0) & " array_obj_ref_259_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_259_data_0));
          --
        end if; 
        if array_obj_ref_259_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_259_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_298_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_298_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_298_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_298_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_298_word_address_0) & " array_obj_ref_298_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_298_data_0));
          --
        end if; 
        if array_obj_ref_298_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_298_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_317_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_317_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_317_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_317_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_317_word_address_0) & " array_obj_ref_317_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_317_data_0));
          --
        end if; 
        if array_obj_ref_317_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_317_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_336_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_336_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_336_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_336_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_336_word_address_0) & " array_obj_ref_336_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_336_data_0));
          --
        end if; 
        if array_obj_ref_336_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_336_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_355_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_355_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_355_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_355_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_355_word_address_0) & " array_obj_ref_355_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_355_data_0));
          --
        end if; 
        if array_obj_ref_355_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_355_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_374_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_374_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_374_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_374_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_374_word_address_0) & " array_obj_ref_374_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_374_data_0));
          --
        end if; 
        if array_obj_ref_374_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_374_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_393_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_393_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_393_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_393_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_393_word_address_0) & " array_obj_ref_393_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_393_data_0));
          --
        end if; 
        if array_obj_ref_393_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_393_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_412_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_412_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_412_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_412_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_412_word_address_0) & " array_obj_ref_412_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_412_data_0));
          --
        end if; 
        if array_obj_ref_412_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_412_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_431_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_431_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_431_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_431_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_431_word_address_0) & " array_obj_ref_431_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_431_data_0));
          --
        end if; 
        if array_obj_ref_431_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_431_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_450_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_450_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_450_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_450_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_450_word_address_0) & " array_obj_ref_450_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_450_data_0));
          --
        end if; 
        if array_obj_ref_450_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_450_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_555_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_555_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_store_0:started:   inputs: " & " array_obj_ref_555_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_555_word_address_0) & " array_obj_ref_555_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_555_data_0));
          --
        end if; 
        if array_obj_ref_555_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_555_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_512_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_512_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_store_0:started:   inputs: " & " array_obj_ref_512_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_512_word_address_0) & " array_obj_ref_512_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_512_data_0));
          --
        end if; 
        if array_obj_ref_512_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_512_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_285_store_0_req_0,
      array_obj_ref_285_store_0_ack_0,
      array_obj_ref_285_store_0_req_1,
      array_obj_ref_285_store_0_ack_1,
      "array_obj_ref_285_store_0",
      "memory_space_1" ,
      array_obj_ref_285_data_0,
      array_obj_ref_285_word_address_0,
      "array_obj_ref_285_data_0",
      "array_obj_ref_285_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_539_store_0_req_0,
      array_obj_ref_539_store_0_ack_0,
      array_obj_ref_539_store_0_req_1,
      array_obj_ref_539_store_0_ack_1,
      "array_obj_ref_539_store_0",
      "memory_space_1" ,
      array_obj_ref_539_data_0,
      array_obj_ref_539_word_address_0,
      "array_obj_ref_539_data_0",
      "array_obj_ref_539_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_272_store_0_req_0,
      array_obj_ref_272_store_0_ack_0,
      array_obj_ref_272_store_0_req_1,
      array_obj_ref_272_store_0_ack_1,
      "array_obj_ref_272_store_0",
      "memory_space_1" ,
      array_obj_ref_272_data_0,
      array_obj_ref_272_word_address_0,
      "array_obj_ref_272_data_0",
      "array_obj_ref_272_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_523_store_0_req_0,
      array_obj_ref_523_store_0_ack_0,
      array_obj_ref_523_store_0_req_1,
      array_obj_ref_523_store_0_ack_1,
      "array_obj_ref_523_store_0",
      "memory_space_1" ,
      array_obj_ref_523_data_0,
      array_obj_ref_523_word_address_0,
      "array_obj_ref_523_data_0",
      "array_obj_ref_523_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_259_store_0_req_0,
      array_obj_ref_259_store_0_ack_0,
      array_obj_ref_259_store_0_req_1,
      array_obj_ref_259_store_0_ack_1,
      "array_obj_ref_259_store_0",
      "memory_space_1" ,
      array_obj_ref_259_data_0,
      array_obj_ref_259_word_address_0,
      "array_obj_ref_259_data_0",
      "array_obj_ref_259_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_298_store_0_req_0,
      array_obj_ref_298_store_0_ack_0,
      array_obj_ref_298_store_0_req_1,
      array_obj_ref_298_store_0_ack_1,
      "array_obj_ref_298_store_0",
      "memory_space_1" ,
      array_obj_ref_298_data_0,
      array_obj_ref_298_word_address_0,
      "array_obj_ref_298_data_0",
      "array_obj_ref_298_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_317_store_0_req_0,
      array_obj_ref_317_store_0_ack_0,
      array_obj_ref_317_store_0_req_1,
      array_obj_ref_317_store_0_ack_1,
      "array_obj_ref_317_store_0",
      "memory_space_1" ,
      array_obj_ref_317_data_0,
      array_obj_ref_317_word_address_0,
      "array_obj_ref_317_data_0",
      "array_obj_ref_317_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_336_store_0_req_0,
      array_obj_ref_336_store_0_ack_0,
      array_obj_ref_336_store_0_req_1,
      array_obj_ref_336_store_0_ack_1,
      "array_obj_ref_336_store_0",
      "memory_space_1" ,
      array_obj_ref_336_data_0,
      array_obj_ref_336_word_address_0,
      "array_obj_ref_336_data_0",
      "array_obj_ref_336_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_355_store_0_req_0,
      array_obj_ref_355_store_0_ack_0,
      array_obj_ref_355_store_0_req_1,
      array_obj_ref_355_store_0_ack_1,
      "array_obj_ref_355_store_0",
      "memory_space_1" ,
      array_obj_ref_355_data_0,
      array_obj_ref_355_word_address_0,
      "array_obj_ref_355_data_0",
      "array_obj_ref_355_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_374_store_0_req_0,
      array_obj_ref_374_store_0_ack_0,
      array_obj_ref_374_store_0_req_1,
      array_obj_ref_374_store_0_ack_1,
      "array_obj_ref_374_store_0",
      "memory_space_1" ,
      array_obj_ref_374_data_0,
      array_obj_ref_374_word_address_0,
      "array_obj_ref_374_data_0",
      "array_obj_ref_374_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_393_store_0_req_0,
      array_obj_ref_393_store_0_ack_0,
      array_obj_ref_393_store_0_req_1,
      array_obj_ref_393_store_0_ack_1,
      "array_obj_ref_393_store_0",
      "memory_space_1" ,
      array_obj_ref_393_data_0,
      array_obj_ref_393_word_address_0,
      "array_obj_ref_393_data_0",
      "array_obj_ref_393_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_412_store_0_req_0,
      array_obj_ref_412_store_0_ack_0,
      array_obj_ref_412_store_0_req_1,
      array_obj_ref_412_store_0_ack_1,
      "array_obj_ref_412_store_0",
      "memory_space_1" ,
      array_obj_ref_412_data_0,
      array_obj_ref_412_word_address_0,
      "array_obj_ref_412_data_0",
      "array_obj_ref_412_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_431_store_0_req_0,
      array_obj_ref_431_store_0_ack_0,
      array_obj_ref_431_store_0_req_1,
      array_obj_ref_431_store_0_ack_1,
      "array_obj_ref_431_store_0",
      "memory_space_1" ,
      array_obj_ref_431_data_0,
      array_obj_ref_431_word_address_0,
      "array_obj_ref_431_data_0",
      "array_obj_ref_431_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_450_store_0_req_0,
      array_obj_ref_450_store_0_ack_0,
      array_obj_ref_450_store_0_req_1,
      array_obj_ref_450_store_0_ack_1,
      "array_obj_ref_450_store_0",
      "memory_space_1" ,
      array_obj_ref_450_data_0,
      array_obj_ref_450_word_address_0,
      "array_obj_ref_450_data_0",
      "array_obj_ref_450_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_555_store_0_req_0,
      array_obj_ref_555_store_0_ack_0,
      array_obj_ref_555_store_0_req_1,
      array_obj_ref_555_store_0_ack_1,
      "array_obj_ref_555_store_0",
      "memory_space_1" ,
      array_obj_ref_555_data_0,
      array_obj_ref_555_word_address_0,
      "array_obj_ref_555_data_0",
      "array_obj_ref_555_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_512_store_0_req_0,
      array_obj_ref_512_store_0_ack_0,
      array_obj_ref_512_store_0_req_1,
      array_obj_ref_512_store_0_ack_1,
      "array_obj_ref_512_store_0",
      "memory_space_1" ,
      array_obj_ref_512_data_0,
      array_obj_ref_512_word_address_0,
      "array_obj_ref_512_data_0",
      "array_obj_ref_512_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_285_store_0 array_obj_ref_539_store_0 array_obj_ref_272_store_0 array_obj_ref_523_store_0 array_obj_ref_259_store_0 array_obj_ref_298_store_0 array_obj_ref_317_store_0 array_obj_ref_336_store_0 array_obj_ref_355_store_0 array_obj_ref_374_store_0 array_obj_ref_393_store_0 array_obj_ref_412_store_0 array_obj_ref_431_store_0 array_obj_ref_450_store_0 array_obj_ref_555_store_0 array_obj_ref_512_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(63 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => true, 3 => true, 4 => true, 5 => true, 6 => true, 7 => true, 8 => true, 9 => true, 10 => true, 11 => true, 12 => false, 13 => true, 14 => false, 15 => true);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= array_obj_ref_285_store_0_req_0;
      reqL_unguarded(14) <= array_obj_ref_539_store_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_272_store_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_523_store_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_259_store_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_298_store_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_317_store_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_336_store_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_355_store_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_374_store_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_393_store_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_412_store_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_431_store_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_450_store_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_555_store_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_512_store_0_req_0;
      array_obj_ref_285_store_0_ack_0 <= ackL_unguarded(15);
      array_obj_ref_539_store_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_272_store_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_523_store_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_259_store_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_298_store_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_317_store_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_336_store_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_355_store_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_374_store_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_393_store_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_412_store_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_431_store_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_450_store_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_555_store_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_512_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= array_obj_ref_285_store_0_req_1;
      reqR_unguarded(14) <= array_obj_ref_539_store_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_272_store_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_523_store_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_259_store_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_298_store_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_317_store_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_336_store_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_355_store_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_374_store_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_393_store_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_412_store_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_431_store_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_450_store_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_555_store_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_512_store_0_req_1;
      array_obj_ref_285_store_0_ack_1 <= ackR_unguarded(15);
      array_obj_ref_539_store_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_272_store_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_523_store_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_259_store_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_298_store_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_317_store_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_336_store_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_355_store_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_374_store_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_393_store_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_412_store_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_431_store_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_450_store_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_555_store_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_512_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  not checkJZero_208(0);
      guard_vector(3)  <=  not checkJZero_208(0);
      guard_vector(4)  <=  not checkJZero_208(0);
      guard_vector(5)  <=  not checkJZero_208(0);
      guard_vector(6)  <=  not checkJZero_208(0);
      guard_vector(7)  <=  not checkJZero_208(0);
      guard_vector(8)  <=  not checkJZero_208(0);
      guard_vector(9)  <=  not checkJZero_208(0);
      guard_vector(10)  <=  not checkJZero_208(0);
      guard_vector(11)  <=  not checkJZero_208(0);
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  not checkJZero_208(0);
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  not checkJZero_208(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_285_word_address_0 & array_obj_ref_539_word_address_0 & array_obj_ref_272_word_address_0 & array_obj_ref_523_word_address_0 & array_obj_ref_259_word_address_0 & array_obj_ref_298_word_address_0 & array_obj_ref_317_word_address_0 & array_obj_ref_336_word_address_0 & array_obj_ref_355_word_address_0 & array_obj_ref_374_word_address_0 & array_obj_ref_393_word_address_0 & array_obj_ref_412_word_address_0 & array_obj_ref_431_word_address_0 & array_obj_ref_450_word_address_0 & array_obj_ref_555_word_address_0 & array_obj_ref_512_word_address_0;
      data_in <= array_obj_ref_285_data_0 & array_obj_ref_539_data_0 & array_obj_ref_272_data_0 & array_obj_ref_523_data_0 & array_obj_ref_259_data_0 & array_obj_ref_298_data_0 & array_obj_ref_317_data_0 & array_obj_ref_336_data_0 & array_obj_ref_355_data_0 & array_obj_ref_374_data_0 & array_obj_ref_393_data_0 & array_obj_ref_412_data_0 & array_obj_ref_431_data_0 & array_obj_ref_450_data_0 & array_obj_ref_555_data_0 & array_obj_ref_512_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(15 downto 0),
          mtag => memory_space_1_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logger for split-operator array_obj_ref_528_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_528_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_store_0:started:   inputs: " & " array_obj_ref_528_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_528_word_address_0) & " array_obj_ref_528_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_528_data_0));
          --
        end if; 
        if array_obj_ref_528_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_528_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_304_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_304_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_304_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_304_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_304_word_address_0) & " array_obj_ref_304_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_304_data_0));
          --
        end if; 
        if array_obj_ref_304_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_304_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_571_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_571_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_store_0:started:   inputs: " & " array_obj_ref_571_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_571_word_address_0) & " array_obj_ref_571_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_571_data_0));
          --
        end if; 
        if array_obj_ref_571_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_571_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_323_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_323_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_323_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_323_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_323_word_address_0) & " array_obj_ref_323_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_323_data_0));
          --
        end if; 
        if array_obj_ref_323_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_323_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_342_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_342_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_342_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_342_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_342_word_address_0) & " array_obj_ref_342_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_342_data_0));
          --
        end if; 
        if array_obj_ref_342_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_342_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_361_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_361_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_361_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_361_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_361_word_address_0) & " array_obj_ref_361_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_361_data_0));
          --
        end if; 
        if array_obj_ref_361_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_361_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_380_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_380_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_380_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_380_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_380_word_address_0) & " array_obj_ref_380_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_380_data_0));
          --
        end if; 
        if array_obj_ref_380_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_380_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_560_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_560_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_store_0:started:   inputs: " & " array_obj_ref_560_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_560_word_address_0) & " array_obj_ref_560_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_560_data_0));
          --
        end if; 
        if array_obj_ref_560_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_560_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_399_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_399_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_399_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_399_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_399_word_address_0) & " array_obj_ref_399_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_399_data_0));
          --
        end if; 
        if array_obj_ref_399_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_399_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_418_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_418_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_418_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_418_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_418_word_address_0) & " array_obj_ref_418_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_418_data_0));
          --
        end if; 
        if array_obj_ref_418_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_418_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_437_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_437_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_437_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_437_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_437_word_address_0) & " array_obj_ref_437_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_437_data_0));
          --
        end if; 
        if array_obj_ref_437_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_437_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_456_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_456_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_456_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_456_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_456_word_address_0) & " array_obj_ref_456_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_456_data_0));
          --
        end if; 
        if array_obj_ref_456_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_456_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_469_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_469_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_469_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_469_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_469_word_address_0) & " array_obj_ref_469_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_469_data_0));
          --
        end if; 
        if array_obj_ref_469_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_469_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_482_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_482_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_482_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_482_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_482_word_address_0) & " array_obj_ref_482_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_482_data_0));
          --
        end if; 
        if array_obj_ref_482_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_482_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_544_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_544_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_store_0:started:   inputs: " & " array_obj_ref_544_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_544_word_address_0) & " array_obj_ref_544_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_544_data_0));
          --
        end if; 
        if array_obj_ref_544_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_544_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_495_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_495_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_495_store_0:started:   inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " array_obj_ref_495_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_495_word_address_0) & " array_obj_ref_495_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_495_data_0));
          --
        end if; 
        if array_obj_ref_495_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:array_obj_ref_495_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_528_store_0_req_0,
      array_obj_ref_528_store_0_ack_0,
      array_obj_ref_528_store_0_req_1,
      array_obj_ref_528_store_0_ack_1,
      "array_obj_ref_528_store_0",
      "memory_space_2" ,
      array_obj_ref_528_data_0,
      array_obj_ref_528_word_address_0,
      "array_obj_ref_528_data_0",
      "array_obj_ref_528_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_304_store_0_req_0,
      array_obj_ref_304_store_0_ack_0,
      array_obj_ref_304_store_0_req_1,
      array_obj_ref_304_store_0_ack_1,
      "array_obj_ref_304_store_0",
      "memory_space_2" ,
      array_obj_ref_304_data_0,
      array_obj_ref_304_word_address_0,
      "array_obj_ref_304_data_0",
      "array_obj_ref_304_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_571_store_0_req_0,
      array_obj_ref_571_store_0_ack_0,
      array_obj_ref_571_store_0_req_1,
      array_obj_ref_571_store_0_ack_1,
      "array_obj_ref_571_store_0",
      "memory_space_2" ,
      array_obj_ref_571_data_0,
      array_obj_ref_571_word_address_0,
      "array_obj_ref_571_data_0",
      "array_obj_ref_571_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_323_store_0_req_0,
      array_obj_ref_323_store_0_ack_0,
      array_obj_ref_323_store_0_req_1,
      array_obj_ref_323_store_0_ack_1,
      "array_obj_ref_323_store_0",
      "memory_space_2" ,
      array_obj_ref_323_data_0,
      array_obj_ref_323_word_address_0,
      "array_obj_ref_323_data_0",
      "array_obj_ref_323_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_342_store_0_req_0,
      array_obj_ref_342_store_0_ack_0,
      array_obj_ref_342_store_0_req_1,
      array_obj_ref_342_store_0_ack_1,
      "array_obj_ref_342_store_0",
      "memory_space_2" ,
      array_obj_ref_342_data_0,
      array_obj_ref_342_word_address_0,
      "array_obj_ref_342_data_0",
      "array_obj_ref_342_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_361_store_0_req_0,
      array_obj_ref_361_store_0_ack_0,
      array_obj_ref_361_store_0_req_1,
      array_obj_ref_361_store_0_ack_1,
      "array_obj_ref_361_store_0",
      "memory_space_2" ,
      array_obj_ref_361_data_0,
      array_obj_ref_361_word_address_0,
      "array_obj_ref_361_data_0",
      "array_obj_ref_361_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_380_store_0_req_0,
      array_obj_ref_380_store_0_ack_0,
      array_obj_ref_380_store_0_req_1,
      array_obj_ref_380_store_0_ack_1,
      "array_obj_ref_380_store_0",
      "memory_space_2" ,
      array_obj_ref_380_data_0,
      array_obj_ref_380_word_address_0,
      "array_obj_ref_380_data_0",
      "array_obj_ref_380_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_560_store_0_req_0,
      array_obj_ref_560_store_0_ack_0,
      array_obj_ref_560_store_0_req_1,
      array_obj_ref_560_store_0_ack_1,
      "array_obj_ref_560_store_0",
      "memory_space_2" ,
      array_obj_ref_560_data_0,
      array_obj_ref_560_word_address_0,
      "array_obj_ref_560_data_0",
      "array_obj_ref_560_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_399_store_0_req_0,
      array_obj_ref_399_store_0_ack_0,
      array_obj_ref_399_store_0_req_1,
      array_obj_ref_399_store_0_ack_1,
      "array_obj_ref_399_store_0",
      "memory_space_2" ,
      array_obj_ref_399_data_0,
      array_obj_ref_399_word_address_0,
      "array_obj_ref_399_data_0",
      "array_obj_ref_399_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_418_store_0_req_0,
      array_obj_ref_418_store_0_ack_0,
      array_obj_ref_418_store_0_req_1,
      array_obj_ref_418_store_0_ack_1,
      "array_obj_ref_418_store_0",
      "memory_space_2" ,
      array_obj_ref_418_data_0,
      array_obj_ref_418_word_address_0,
      "array_obj_ref_418_data_0",
      "array_obj_ref_418_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_437_store_0_req_0,
      array_obj_ref_437_store_0_ack_0,
      array_obj_ref_437_store_0_req_1,
      array_obj_ref_437_store_0_ack_1,
      "array_obj_ref_437_store_0",
      "memory_space_2" ,
      array_obj_ref_437_data_0,
      array_obj_ref_437_word_address_0,
      "array_obj_ref_437_data_0",
      "array_obj_ref_437_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_456_store_0_req_0,
      array_obj_ref_456_store_0_ack_0,
      array_obj_ref_456_store_0_req_1,
      array_obj_ref_456_store_0_ack_1,
      "array_obj_ref_456_store_0",
      "memory_space_2" ,
      array_obj_ref_456_data_0,
      array_obj_ref_456_word_address_0,
      "array_obj_ref_456_data_0",
      "array_obj_ref_456_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_469_store_0_req_0,
      array_obj_ref_469_store_0_ack_0,
      array_obj_ref_469_store_0_req_1,
      array_obj_ref_469_store_0_ack_1,
      "array_obj_ref_469_store_0",
      "memory_space_2" ,
      array_obj_ref_469_data_0,
      array_obj_ref_469_word_address_0,
      "array_obj_ref_469_data_0",
      "array_obj_ref_469_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_482_store_0_req_0,
      array_obj_ref_482_store_0_ack_0,
      array_obj_ref_482_store_0_req_1,
      array_obj_ref_482_store_0_ack_1,
      "array_obj_ref_482_store_0",
      "memory_space_2" ,
      array_obj_ref_482_data_0,
      array_obj_ref_482_word_address_0,
      "array_obj_ref_482_data_0",
      "array_obj_ref_482_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_544_store_0_req_0,
      array_obj_ref_544_store_0_ack_0,
      array_obj_ref_544_store_0_req_1,
      array_obj_ref_544_store_0_ack_1,
      "array_obj_ref_544_store_0",
      "memory_space_2" ,
      array_obj_ref_544_data_0,
      array_obj_ref_544_word_address_0,
      "array_obj_ref_544_data_0",
      "array_obj_ref_544_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_495_store_0_req_0,
      array_obj_ref_495_store_0_ack_0,
      array_obj_ref_495_store_0_req_1,
      array_obj_ref_495_store_0_ack_1,
      "array_obj_ref_495_store_0",
      "memory_space_2" ,
      array_obj_ref_495_data_0,
      array_obj_ref_495_word_address_0,
      "array_obj_ref_495_data_0",
      "array_obj_ref_495_word_address_0" -- 
    );
    -- shared store operator group (1) : array_obj_ref_528_store_0 array_obj_ref_304_store_0 array_obj_ref_571_store_0 array_obj_ref_323_store_0 array_obj_ref_342_store_0 array_obj_ref_361_store_0 array_obj_ref_380_store_0 array_obj_ref_560_store_0 array_obj_ref_399_store_0 array_obj_ref_418_store_0 array_obj_ref_437_store_0 array_obj_ref_456_store_0 array_obj_ref_469_store_0 array_obj_ref_482_store_0 array_obj_ref_544_store_0 array_obj_ref_495_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(63 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => true, 1 => false, 2 => true, 3 => true, 4 => true, 5 => true, 6 => true, 7 => true, 8 => false, 9 => true, 10 => true, 11 => true, 12 => true, 13 => false, 14 => true, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= array_obj_ref_528_store_0_req_0;
      reqL_unguarded(14) <= array_obj_ref_304_store_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_571_store_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_323_store_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_342_store_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_361_store_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_380_store_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_560_store_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_399_store_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_418_store_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_437_store_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_456_store_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_469_store_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_482_store_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_544_store_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_495_store_0_req_0;
      array_obj_ref_528_store_0_ack_0 <= ackL_unguarded(15);
      array_obj_ref_304_store_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_571_store_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_323_store_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_342_store_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_361_store_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_380_store_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_560_store_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_399_store_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_418_store_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_437_store_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_456_store_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_469_store_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_482_store_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_544_store_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_495_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= array_obj_ref_528_store_0_req_1;
      reqR_unguarded(14) <= array_obj_ref_304_store_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_571_store_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_323_store_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_342_store_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_361_store_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_380_store_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_560_store_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_399_store_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_418_store_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_437_store_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_456_store_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_469_store_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_482_store_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_544_store_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_495_store_0_req_1;
      array_obj_ref_528_store_0_ack_1 <= ackR_unguarded(15);
      array_obj_ref_304_store_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_571_store_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_323_store_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_342_store_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_361_store_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_380_store_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_560_store_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_399_store_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_418_store_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_437_store_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_456_store_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_469_store_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_482_store_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_544_store_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_495_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not checkJZero_208(0);
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  not checkJZero_208(0);
      guard_vector(3)  <=  not checkJZero_208(0);
      guard_vector(4)  <=  not checkJZero_208(0);
      guard_vector(5)  <=  not checkJZero_208(0);
      guard_vector(6)  <=  not checkJZero_208(0);
      guard_vector(7)  <=  not checkJZero_208(0);
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  not checkJZero_208(0);
      guard_vector(10)  <=  not checkJZero_208(0);
      guard_vector(11)  <=  not checkJZero_208(0);
      guard_vector(12)  <=  not checkJZero_208(0);
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  not checkJZero_208(0);
      guard_vector(15)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_528_word_address_0 & array_obj_ref_304_word_address_0 & array_obj_ref_571_word_address_0 & array_obj_ref_323_word_address_0 & array_obj_ref_342_word_address_0 & array_obj_ref_361_word_address_0 & array_obj_ref_380_word_address_0 & array_obj_ref_560_word_address_0 & array_obj_ref_399_word_address_0 & array_obj_ref_418_word_address_0 & array_obj_ref_437_word_address_0 & array_obj_ref_456_word_address_0 & array_obj_ref_469_word_address_0 & array_obj_ref_482_word_address_0 & array_obj_ref_544_word_address_0 & array_obj_ref_495_word_address_0;
      data_in <= array_obj_ref_528_data_0 & array_obj_ref_304_data_0 & array_obj_ref_571_data_0 & array_obj_ref_323_data_0 & array_obj_ref_342_data_0 & array_obj_ref_361_data_0 & array_obj_ref_380_data_0 & array_obj_ref_560_data_0 & array_obj_ref_399_data_0 & array_obj_ref_418_data_0 & array_obj_ref_437_data_0 & array_obj_ref_456_data_0 & array_obj_ref_469_data_0 & array_obj_ref_482_data_0 & array_obj_ref_544_data_0 & array_obj_ref_495_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 4,
        data_width => 16,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(3 downto 0),
          mdata => memory_space_2_sr_data(15 downto 0),
          mtag => memory_space_2_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- logger for split-operator call_stmt_281_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_281_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_281_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_276_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_276_wire_constant) & " rowI_212 = "& Convert_SLV_To_Hex_String(rowI_212) & " col2_248 = "& Convert_SLV_To_Hex_String(col2_248) & " R_write_data_zero_279_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_279_wire_constant));
          --
        end if; 
        if call_stmt_281_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_281_call:finished:  outputs: " & " rdata_I02_281= "  & Convert_SLV_To_Hex_String(rdata_I02_281));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_294_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_294_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_294_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_289_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_289_wire_constant) & " rowI_1_218 = "& Convert_SLV_To_Hex_String(rowI_1_218) & " col0_240 = "& Convert_SLV_To_Hex_String(col0_240) & " R_write_data_zero_292_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_292_wire_constant));
          --
        end if; 
        if call_stmt_294_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_294_call:finished:  outputs: " & " rdata_I10_294= "  & Convert_SLV_To_Hex_String(rdata_I10_294));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_255_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_255_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_255_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_250_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_250_wire_constant) & " rowI_212 = "& Convert_SLV_To_Hex_String(rowI_212) & " col0_240 = "& Convert_SLV_To_Hex_String(col0_240) & " R_write_data_zero_253_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_253_wire_constant));
          --
        end if; 
        if call_stmt_255_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_255_call:finished:  outputs: " & " rdata_I00_255= "  & Convert_SLV_To_Hex_String(rdata_I00_255));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_536_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_536_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_536_call:started:  Call to module accessMem inputs: " & " R_read_signal_531_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_531_wire_constant) & " rowI_2_224 = "& Convert_SLV_To_Hex_String(rowI_2_224) & " J_3_503 = "& Convert_SLV_To_Hex_String(J_3_503) & " R_write_data_zero_534_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_534_wire_constant));
          --
        end if; 
        if call_stmt_536_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_536_call:finished:  outputs: " & " rdata_ifmap2_536= "  & Convert_SLV_To_Hex_String(rdata_ifmap2_536));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_268_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_268_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_268_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_263_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_263_wire_constant) & " rowI_212 = "& Convert_SLV_To_Hex_String(rowI_212) & " col1_244 = "& Convert_SLV_To_Hex_String(col1_244) & " R_write_data_zero_266_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_266_wire_constant));
          --
        end if; 
        if call_stmt_268_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_268_call:finished:  outputs: " & " rdata_I01_268= "  & Convert_SLV_To_Hex_String(rdata_I01_268));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_552_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_552_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_552_call:started:  Call to module accessMem inputs: " & " R_read_signal_547_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_547_wire_constant) & " rowI_3_230 = "& Convert_SLV_To_Hex_String(rowI_3_230) & " J_3_503 = "& Convert_SLV_To_Hex_String(J_3_503) & " R_write_data_zero_550_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_550_wire_constant));
          --
        end if; 
        if call_stmt_552_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_552_call:finished:  outputs: " & " rdata_ifmap3_552= "  & Convert_SLV_To_Hex_String(rdata_ifmap3_552));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_313_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_313_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_313_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_308_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_308_wire_constant) & " rowI_1_218 = "& Convert_SLV_To_Hex_String(rowI_1_218) & " col1_244 = "& Convert_SLV_To_Hex_String(col1_244) & " R_write_data_zero_311_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_311_wire_constant));
          --
        end if; 
        if call_stmt_313_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_313_call:finished:  outputs: " & " rdata_I11_313= "  & Convert_SLV_To_Hex_String(rdata_I11_313));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_332_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_332_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_332_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_327_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_327_wire_constant) & " rowI_1_218 = "& Convert_SLV_To_Hex_String(rowI_1_218) & " col2_248 = "& Convert_SLV_To_Hex_String(col2_248) & " R_write_data_zero_330_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_330_wire_constant));
          --
        end if; 
        if call_stmt_332_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_332_call:finished:  outputs: " & " rdata_I12_332= "  & Convert_SLV_To_Hex_String(rdata_I12_332));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_351_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_351_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_351_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_346_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_346_wire_constant) & " rowI_2_224 = "& Convert_SLV_To_Hex_String(rowI_2_224) & " col0_240 = "& Convert_SLV_To_Hex_String(col0_240) & " R_write_data_zero_349_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_349_wire_constant));
          --
        end if; 
        if call_stmt_351_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_351_call:finished:  outputs: " & " rdata_I20_351= "  & Convert_SLV_To_Hex_String(rdata_I20_351));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_370_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_370_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_370_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_365_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_365_wire_constant) & " rowI_2_224 = "& Convert_SLV_To_Hex_String(rowI_2_224) & " col1_244 = "& Convert_SLV_To_Hex_String(col1_244) & " R_write_data_zero_368_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_368_wire_constant));
          --
        end if; 
        if call_stmt_370_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_370_call:finished:  outputs: " & " rdata_I21_370= "  & Convert_SLV_To_Hex_String(rdata_I21_370));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_568_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_568_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_568_call:started:  Call to module accessMem inputs: " & " R_read_signal_563_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_563_wire_constant) & " rowI_4_236 = "& Convert_SLV_To_Hex_String(rowI_4_236) & " J_3_503 = "& Convert_SLV_To_Hex_String(J_3_503) & " R_write_data_zero_566_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_566_wire_constant));
          --
        end if; 
        if call_stmt_568_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_568_call:finished:  outputs: " & " rdata_ifmap4_568= "  & Convert_SLV_To_Hex_String(rdata_ifmap4_568));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_389_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_389_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_389_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_384_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_384_wire_constant) & " rowI_2_224 = "& Convert_SLV_To_Hex_String(rowI_2_224) & " col2_248 = "& Convert_SLV_To_Hex_String(col2_248) & " R_write_data_zero_387_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_387_wire_constant));
          --
        end if; 
        if call_stmt_389_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_389_call:finished:  outputs: " & " rdata_I22_389= "  & Convert_SLV_To_Hex_String(rdata_I22_389));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_408_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_408_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_408_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_403_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_403_wire_constant) & " rowI_3_230 = "& Convert_SLV_To_Hex_String(rowI_3_230) & " col0_240 = "& Convert_SLV_To_Hex_String(col0_240) & " R_write_data_zero_406_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_406_wire_constant));
          --
        end if; 
        if call_stmt_408_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_408_call:finished:  outputs: " & " rdata_I30_408= "  & Convert_SLV_To_Hex_String(rdata_I30_408));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_427_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_427_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_427_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_422_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_422_wire_constant) & " rowI_3_230 = "& Convert_SLV_To_Hex_String(rowI_3_230) & " col1_244 = "& Convert_SLV_To_Hex_String(col1_244) & " R_write_data_zero_425_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_425_wire_constant));
          --
        end if; 
        if call_stmt_427_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_427_call:finished:  outputs: " & " rdata_I31_427= "  & Convert_SLV_To_Hex_String(rdata_I31_427));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_446_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_446_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_446_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_441_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_441_wire_constant) & " rowI_3_230 = "& Convert_SLV_To_Hex_String(rowI_3_230) & " col2_248 = "& Convert_SLV_To_Hex_String(col2_248) & " R_write_data_zero_444_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_444_wire_constant));
          --
        end if; 
        if call_stmt_446_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_446_call:finished:  outputs: " & " rdata_I32_446= "  & Convert_SLV_To_Hex_String(rdata_I32_446));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_465_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_465_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_465_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_460_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_460_wire_constant) & " rowI_4_236 = "& Convert_SLV_To_Hex_String(rowI_4_236) & " col0_240 = "& Convert_SLV_To_Hex_String(col0_240) & " R_write_data_zero_463_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_463_wire_constant));
          --
        end if; 
        if call_stmt_465_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_465_call:finished:  outputs: " & " rdata_I40_465= "  & Convert_SLV_To_Hex_String(rdata_I40_465));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_478_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_478_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_478_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_473_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_473_wire_constant) & " rowI_4_236 = "& Convert_SLV_To_Hex_String(rowI_4_236) & " col1_244 = "& Convert_SLV_To_Hex_String(col1_244) & " R_write_data_zero_476_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_476_wire_constant));
          --
        end if; 
        if call_stmt_478_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_478_call:finished:  outputs: " & " rdata_I41_478= "  & Convert_SLV_To_Hex_String(rdata_I41_478));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_491_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_491_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_491_call:started:  Call to module accessMem inputs: " & " checkJZero_208 (guard complement )= " & Convert_SLV_To_String(checkJZero_208) & " R_read_signal_486_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_486_wire_constant) & " rowI_4_236 = "& Convert_SLV_To_Hex_String(rowI_4_236) & " col2_248 = "& Convert_SLV_To_Hex_String(col2_248) & " R_write_data_zero_489_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_489_wire_constant));
          --
        end if; 
        if call_stmt_491_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_491_call:finished:  outputs: " & " rdata_I42_491= "  & Convert_SLV_To_Hex_String(rdata_I42_491));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_509_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_509_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_509_call:started:  Call to module accessMem inputs: " & " R_read_signal_504_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_504_wire_constant) & " rowI_212 = "& Convert_SLV_To_Hex_String(rowI_212) & " J_3_503 = "& Convert_SLV_To_Hex_String(J_3_503) & " R_write_data_zero_507_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_507_wire_constant));
          --
        end if; 
        if call_stmt_509_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_509_call:finished:  outputs: " & " rdata_ifmap0_509= "  & Convert_SLV_To_Hex_String(rdata_ifmap0_509));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_520_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_520_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_520_call:started:  Call to module accessMem inputs: " & " R_read_signal_515_wire_constant = "& Convert_SLV_To_Hex_String(R_read_signal_515_wire_constant) & " rowI_1_218 = "& Convert_SLV_To_Hex_String(rowI_1_218) & " J_3_503 = "& Convert_SLV_To_Hex_String(J_3_503) & " R_write_data_zero_518_wire_constant = "& Convert_SLV_To_Hex_String(R_write_data_zero_518_wire_constant));
          --
        end if; 
        if call_stmt_520_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:initIfMaps:DP:call_stmt_520_call:finished:  outputs: " & " rdata_ifmap1_520= "  & Convert_SLV_To_Hex_String(rdata_ifmap1_520));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_281_call call_stmt_294_call call_stmt_255_call call_stmt_536_call call_stmt_268_call call_stmt_552_call call_stmt_313_call call_stmt_332_call call_stmt_351_call call_stmt_370_call call_stmt_568_call call_stmt_389_call call_stmt_408_call call_stmt_427_call call_stmt_446_call call_stmt_465_call call_stmt_478_call call_stmt_491_call call_stmt_509_call call_stmt_520_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(559 downto 0);
      signal data_out: std_logic_vector(319 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 19 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 19 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 19 downto 0);
      signal guard_vector : std_logic_vector( 19 downto 0);
      constant inBUFs : IntegerArray(19 downto 0) := (19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(19 downto 0) := (19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(19 downto 0) := (0 => false, 1 => false, 2 => true, 3 => true, 4 => true, 5 => true, 6 => true, 7 => true, 8 => true, 9 => false, 10 => true, 11 => true, 12 => true, 13 => true, 14 => false, 15 => true, 16 => false, 17 => true, 18 => true, 19 => true);
      constant guardBuffering: IntegerArray(19 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2);
      -- 
    begin -- 
      reqL_unguarded(19) <= call_stmt_281_call_req_0;
      reqL_unguarded(18) <= call_stmt_294_call_req_0;
      reqL_unguarded(17) <= call_stmt_255_call_req_0;
      reqL_unguarded(16) <= call_stmt_536_call_req_0;
      reqL_unguarded(15) <= call_stmt_268_call_req_0;
      reqL_unguarded(14) <= call_stmt_552_call_req_0;
      reqL_unguarded(13) <= call_stmt_313_call_req_0;
      reqL_unguarded(12) <= call_stmt_332_call_req_0;
      reqL_unguarded(11) <= call_stmt_351_call_req_0;
      reqL_unguarded(10) <= call_stmt_370_call_req_0;
      reqL_unguarded(9) <= call_stmt_568_call_req_0;
      reqL_unguarded(8) <= call_stmt_389_call_req_0;
      reqL_unguarded(7) <= call_stmt_408_call_req_0;
      reqL_unguarded(6) <= call_stmt_427_call_req_0;
      reqL_unguarded(5) <= call_stmt_446_call_req_0;
      reqL_unguarded(4) <= call_stmt_465_call_req_0;
      reqL_unguarded(3) <= call_stmt_478_call_req_0;
      reqL_unguarded(2) <= call_stmt_491_call_req_0;
      reqL_unguarded(1) <= call_stmt_509_call_req_0;
      reqL_unguarded(0) <= call_stmt_520_call_req_0;
      call_stmt_281_call_ack_0 <= ackL_unguarded(19);
      call_stmt_294_call_ack_0 <= ackL_unguarded(18);
      call_stmt_255_call_ack_0 <= ackL_unguarded(17);
      call_stmt_536_call_ack_0 <= ackL_unguarded(16);
      call_stmt_268_call_ack_0 <= ackL_unguarded(15);
      call_stmt_552_call_ack_0 <= ackL_unguarded(14);
      call_stmt_313_call_ack_0 <= ackL_unguarded(13);
      call_stmt_332_call_ack_0 <= ackL_unguarded(12);
      call_stmt_351_call_ack_0 <= ackL_unguarded(11);
      call_stmt_370_call_ack_0 <= ackL_unguarded(10);
      call_stmt_568_call_ack_0 <= ackL_unguarded(9);
      call_stmt_389_call_ack_0 <= ackL_unguarded(8);
      call_stmt_408_call_ack_0 <= ackL_unguarded(7);
      call_stmt_427_call_ack_0 <= ackL_unguarded(6);
      call_stmt_446_call_ack_0 <= ackL_unguarded(5);
      call_stmt_465_call_ack_0 <= ackL_unguarded(4);
      call_stmt_478_call_ack_0 <= ackL_unguarded(3);
      call_stmt_491_call_ack_0 <= ackL_unguarded(2);
      call_stmt_509_call_ack_0 <= ackL_unguarded(1);
      call_stmt_520_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(19) <= call_stmt_281_call_req_1;
      reqR_unguarded(18) <= call_stmt_294_call_req_1;
      reqR_unguarded(17) <= call_stmt_255_call_req_1;
      reqR_unguarded(16) <= call_stmt_536_call_req_1;
      reqR_unguarded(15) <= call_stmt_268_call_req_1;
      reqR_unguarded(14) <= call_stmt_552_call_req_1;
      reqR_unguarded(13) <= call_stmt_313_call_req_1;
      reqR_unguarded(12) <= call_stmt_332_call_req_1;
      reqR_unguarded(11) <= call_stmt_351_call_req_1;
      reqR_unguarded(10) <= call_stmt_370_call_req_1;
      reqR_unguarded(9) <= call_stmt_568_call_req_1;
      reqR_unguarded(8) <= call_stmt_389_call_req_1;
      reqR_unguarded(7) <= call_stmt_408_call_req_1;
      reqR_unguarded(6) <= call_stmt_427_call_req_1;
      reqR_unguarded(5) <= call_stmt_446_call_req_1;
      reqR_unguarded(4) <= call_stmt_465_call_req_1;
      reqR_unguarded(3) <= call_stmt_478_call_req_1;
      reqR_unguarded(2) <= call_stmt_491_call_req_1;
      reqR_unguarded(1) <= call_stmt_509_call_req_1;
      reqR_unguarded(0) <= call_stmt_520_call_req_1;
      call_stmt_281_call_ack_1 <= ackR_unguarded(19);
      call_stmt_294_call_ack_1 <= ackR_unguarded(18);
      call_stmt_255_call_ack_1 <= ackR_unguarded(17);
      call_stmt_536_call_ack_1 <= ackR_unguarded(16);
      call_stmt_268_call_ack_1 <= ackR_unguarded(15);
      call_stmt_552_call_ack_1 <= ackR_unguarded(14);
      call_stmt_313_call_ack_1 <= ackR_unguarded(13);
      call_stmt_332_call_ack_1 <= ackR_unguarded(12);
      call_stmt_351_call_ack_1 <= ackR_unguarded(11);
      call_stmt_370_call_ack_1 <= ackR_unguarded(10);
      call_stmt_568_call_ack_1 <= ackR_unguarded(9);
      call_stmt_389_call_ack_1 <= ackR_unguarded(8);
      call_stmt_408_call_ack_1 <= ackR_unguarded(7);
      call_stmt_427_call_ack_1 <= ackR_unguarded(6);
      call_stmt_446_call_ack_1 <= ackR_unguarded(5);
      call_stmt_465_call_ack_1 <= ackR_unguarded(4);
      call_stmt_478_call_ack_1 <= ackR_unguarded(3);
      call_stmt_491_call_ack_1 <= ackR_unguarded(2);
      call_stmt_509_call_ack_1 <= ackR_unguarded(1);
      call_stmt_520_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  not checkJZero_208(0);
      guard_vector(3)  <=  not checkJZero_208(0);
      guard_vector(4)  <=  not checkJZero_208(0);
      guard_vector(5)  <=  not checkJZero_208(0);
      guard_vector(6)  <=  not checkJZero_208(0);
      guard_vector(7)  <=  not checkJZero_208(0);
      guard_vector(8)  <=  not checkJZero_208(0);
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  not checkJZero_208(0);
      guard_vector(11)  <=  not checkJZero_208(0);
      guard_vector(12)  <=  not checkJZero_208(0);
      guard_vector(13)  <=  not checkJZero_208(0);
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  not checkJZero_208(0);
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  not checkJZero_208(0);
      guard_vector(18)  <=  not checkJZero_208(0);
      guard_vector(19)  <=  not checkJZero_208(0);
      accessMem_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_4: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_5: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_6: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_7: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_8: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_9: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_10: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_11: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_12: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_13: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_14: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_15: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_16: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_16", num_slots => 1) -- 
        port map (req => reqL_unregulated(16), -- 
          ack => ackL_unregulated(16),
          regulated_req => reqL(16),
          regulated_ack => ackL(16),
          release_req => reqR(16),
          release_ack => ackR(16),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_17: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_17", num_slots => 1) -- 
        port map (req => reqL_unregulated(17), -- 
          ack => ackL_unregulated(17),
          regulated_req => reqL(17),
          regulated_ack => ackL(17),
          release_req => reqR(17),
          release_ack => ackR(17),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_18: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_18", num_slots => 1) -- 
        port map (req => reqL_unregulated(18), -- 
          ack => ackL_unregulated(18),
          regulated_req => reqL(18),
          regulated_ack => ackL(18),
          release_req => reqR(18),
          release_ack => ackR(18),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_accessRegulator_19: access_regulator_base generic map (name => "accessMem_call_group_0_accessRegulator_19", num_slots => 1) -- 
        port map (req => reqL_unregulated(19), -- 
          ack => ackL_unregulated(19),
          regulated_req => reqL(19),
          regulated_ack => ackL(19),
          release_req => reqR(19),
          release_ack => ackR(19),
          clk => clk, reset => reset); -- 
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 20, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= R_read_signal_276_wire_constant & rowI_212 & col2_248 & R_write_data_zero_279_wire_constant & R_read_signal_289_wire_constant & rowI_1_218 & col0_240 & R_write_data_zero_292_wire_constant & R_read_signal_250_wire_constant & rowI_212 & col0_240 & R_write_data_zero_253_wire_constant & R_read_signal_531_wire_constant & rowI_2_224 & J_3_503 & R_write_data_zero_534_wire_constant & R_read_signal_263_wire_constant & rowI_212 & col1_244 & R_write_data_zero_266_wire_constant & R_read_signal_547_wire_constant & rowI_3_230 & J_3_503 & R_write_data_zero_550_wire_constant & R_read_signal_308_wire_constant & rowI_1_218 & col1_244 & R_write_data_zero_311_wire_constant & R_read_signal_327_wire_constant & rowI_1_218 & col2_248 & R_write_data_zero_330_wire_constant & R_read_signal_346_wire_constant & rowI_2_224 & col0_240 & R_write_data_zero_349_wire_constant & R_read_signal_365_wire_constant & rowI_2_224 & col1_244 & R_write_data_zero_368_wire_constant & R_read_signal_563_wire_constant & rowI_4_236 & J_3_503 & R_write_data_zero_566_wire_constant & R_read_signal_384_wire_constant & rowI_2_224 & col2_248 & R_write_data_zero_387_wire_constant & R_read_signal_403_wire_constant & rowI_3_230 & col0_240 & R_write_data_zero_406_wire_constant & R_read_signal_422_wire_constant & rowI_3_230 & col1_244 & R_write_data_zero_425_wire_constant & R_read_signal_441_wire_constant & rowI_3_230 & col2_248 & R_write_data_zero_444_wire_constant & R_read_signal_460_wire_constant & rowI_4_236 & col0_240 & R_write_data_zero_463_wire_constant & R_read_signal_473_wire_constant & rowI_4_236 & col1_244 & R_write_data_zero_476_wire_constant & R_read_signal_486_wire_constant & rowI_4_236 & col2_248 & R_write_data_zero_489_wire_constant & R_read_signal_504_wire_constant & rowI_212 & J_3_503 & R_write_data_zero_507_wire_constant & R_read_signal_515_wire_constant & rowI_1_218 & J_3_503 & R_write_data_zero_518_wire_constant;
      rdata_I02_281 <= data_out(319 downto 304);
      rdata_I10_294 <= data_out(303 downto 288);
      rdata_I00_255 <= data_out(287 downto 272);
      rdata_ifmap2_536 <= data_out(271 downto 256);
      rdata_I01_268 <= data_out(255 downto 240);
      rdata_ifmap3_552 <= data_out(239 downto 224);
      rdata_I11_313 <= data_out(223 downto 208);
      rdata_I12_332 <= data_out(207 downto 192);
      rdata_I20_351 <= data_out(191 downto 176);
      rdata_I21_370 <= data_out(175 downto 160);
      rdata_ifmap4_568 <= data_out(159 downto 144);
      rdata_I22_389 <= data_out(143 downto 128);
      rdata_I30_408 <= data_out(127 downto 112);
      rdata_I31_427 <= data_out(111 downto 96);
      rdata_I32_446 <= data_out(95 downto 80);
      rdata_I40_465 <= data_out(79 downto 64);
      rdata_I41_478 <= data_out(63 downto 48);
      rdata_I42_491 <= data_out(47 downto 32);
      rdata_ifmap0_509 <= data_out(31 downto 16);
      rdata_ifmap1_520 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 560,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 5,
        nreqs => 20,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 320,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 20) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end initIfMaps_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity mainAcc is -- 
  generic (tag_length : integer); 
  port ( -- 
    I : in  std_logic_vector(5 downto 0);
    J : in  std_logic_vector(4 downto 0);
    col_to_be_replaced : in  std_logic_vector(1 downto 0);
    ofmap_pixel : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mainAcc;
architecture mainAcc_arch of mainAcc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 13)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal I_buffer :  std_logic_vector(5 downto 0);
  signal I_update_enable: Boolean;
  signal J_buffer :  std_logic_vector(4 downto 0);
  signal J_update_enable: Boolean;
  signal col_to_be_replaced_buffer :  std_logic_vector(1 downto 0);
  signal col_to_be_replaced_update_enable: Boolean;
  -- output port buffer signals
  signal ofmap_pixel_buffer :  std_logic_vector(15 downto 0);
  signal ofmap_pixel_update_enable: Boolean;
  signal mainAcc_CP_2438_start: Boolean;
  signal mainAcc_CP_2438_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_708_load_0_req_0 : boolean;
  signal array_obj_ref_691_load_0_ack_0 : boolean;
  signal array_obj_ref_691_load_0_ack_1 : boolean;
  signal array_obj_ref_691_load_0_req_0 : boolean;
  signal array_obj_ref_691_load_0_req_1 : boolean;
  signal array_obj_ref_688_index_offset_ack_1 : boolean;
  signal type_cast_693_inst_ack_0 : boolean;
  signal array_obj_ref_698_load_0_req_1 : boolean;
  signal type_cast_693_inst_req_0 : boolean;
  signal array_obj_ref_698_index_offset_req_1 : boolean;
  signal array_obj_ref_688_index_offset_ack_0 : boolean;
  signal array_obj_ref_708_index_offset_req_0 : boolean;
  signal array_obj_ref_688_load_0_req_0 : boolean;
  signal type_cast_803_inst_ack_1 : boolean;
  signal array_obj_ref_698_index_offset_ack_1 : boolean;
  signal array_obj_ref_708_index_offset_ack_1 : boolean;
  signal type_cast_703_inst_req_0 : boolean;
  signal type_cast_703_inst_ack_0 : boolean;
  signal array_obj_ref_708_index_offset_ack_0 : boolean;
  signal array_obj_ref_698_load_0_ack_1 : boolean;
  signal type_cast_703_inst_req_1 : boolean;
  signal type_cast_703_inst_ack_1 : boolean;
  signal array_obj_ref_701_load_0_req_1 : boolean;
  signal type_cast_693_inst_ack_1 : boolean;
  signal type_cast_693_inst_req_1 : boolean;
  signal array_obj_ref_798_load_0_req_1 : boolean;
  signal array_obj_ref_688_load_0_ack_0 : boolean;
  signal array_obj_ref_711_load_0_req_0 : boolean;
  signal array_obj_ref_711_load_0_ack_0 : boolean;
  signal array_obj_ref_698_load_0_ack_0 : boolean;
  signal array_obj_ref_708_load_0_req_1 : boolean;
  signal array_obj_ref_688_index_offset_req_0 : boolean;
  signal array_obj_ref_698_index_offset_req_0 : boolean;
  signal array_obj_ref_708_index_offset_req_1 : boolean;
  signal array_obj_ref_701_load_0_ack_1 : boolean;
  signal array_obj_ref_688_index_offset_req_1 : boolean;
  signal array_obj_ref_698_load_0_req_0 : boolean;
  signal array_obj_ref_801_load_0_ack_1 : boolean;
  signal array_obj_ref_698_index_offset_ack_0 : boolean;
  signal array_obj_ref_708_load_0_ack_1 : boolean;
  signal array_obj_ref_701_load_0_ack_0 : boolean;
  signal array_obj_ref_708_load_0_ack_0 : boolean;
  signal array_obj_ref_688_load_0_ack_1 : boolean;
  signal array_obj_ref_701_load_0_req_0 : boolean;
  signal array_obj_ref_688_load_0_req_1 : boolean;
  signal array_obj_ref_801_load_0_req_1 : boolean;
  signal array_obj_ref_711_load_0_ack_1 : boolean;
  signal array_obj_ref_711_load_0_req_1 : boolean;
  signal array_obj_ref_798_load_0_ack_1 : boolean;
  signal type_cast_803_inst_req_0 : boolean;
  signal type_cast_803_inst_ack_0 : boolean;
  signal MUX_647_inst_req_0 : boolean;
  signal MUX_647_inst_ack_0 : boolean;
  signal MUX_647_inst_req_1 : boolean;
  signal MUX_647_inst_ack_1 : boolean;
  signal MUX_661_inst_req_0 : boolean;
  signal MUX_661_inst_ack_0 : boolean;
  signal MUX_661_inst_req_1 : boolean;
  signal MUX_661_inst_ack_1 : boolean;
  signal type_cast_803_inst_req_1 : boolean;
  signal MUX_673_inst_req_0 : boolean;
  signal MUX_673_inst_ack_0 : boolean;
  signal MUX_673_inst_req_1 : boolean;
  signal MUX_673_inst_ack_1 : boolean;
  signal array_obj_ref_678_index_offset_req_0 : boolean;
  signal array_obj_ref_678_index_offset_ack_0 : boolean;
  signal array_obj_ref_678_index_offset_req_1 : boolean;
  signal array_obj_ref_678_index_offset_ack_1 : boolean;
  signal array_obj_ref_678_load_0_req_0 : boolean;
  signal array_obj_ref_678_load_0_ack_0 : boolean;
  signal array_obj_ref_678_load_0_req_1 : boolean;
  signal array_obj_ref_678_load_0_ack_1 : boolean;
  signal array_obj_ref_681_load_0_req_0 : boolean;
  signal array_obj_ref_681_load_0_ack_0 : boolean;
  signal array_obj_ref_681_load_0_req_1 : boolean;
  signal array_obj_ref_681_load_0_ack_1 : boolean;
  signal type_cast_683_inst_req_0 : boolean;
  signal type_cast_683_inst_ack_0 : boolean;
  signal type_cast_683_inst_req_1 : boolean;
  signal type_cast_683_inst_ack_1 : boolean;
  signal type_cast_713_inst_req_0 : boolean;
  signal type_cast_713_inst_ack_0 : boolean;
  signal type_cast_713_inst_req_1 : boolean;
  signal type_cast_713_inst_ack_1 : boolean;
  signal array_obj_ref_718_index_offset_req_0 : boolean;
  signal array_obj_ref_718_index_offset_ack_0 : boolean;
  signal array_obj_ref_718_index_offset_req_1 : boolean;
  signal array_obj_ref_718_index_offset_ack_1 : boolean;
  signal array_obj_ref_718_load_0_req_0 : boolean;
  signal array_obj_ref_718_load_0_ack_0 : boolean;
  signal array_obj_ref_718_load_0_req_1 : boolean;
  signal array_obj_ref_718_load_0_ack_1 : boolean;
  signal array_obj_ref_721_load_0_req_0 : boolean;
  signal array_obj_ref_721_load_0_ack_0 : boolean;
  signal array_obj_ref_721_load_0_req_1 : boolean;
  signal array_obj_ref_721_load_0_ack_1 : boolean;
  signal type_cast_723_inst_req_0 : boolean;
  signal type_cast_723_inst_ack_0 : boolean;
  signal type_cast_723_inst_req_1 : boolean;
  signal type_cast_723_inst_ack_1 : boolean;
  signal array_obj_ref_728_index_offset_req_0 : boolean;
  signal array_obj_ref_728_index_offset_ack_0 : boolean;
  signal array_obj_ref_728_index_offset_req_1 : boolean;
  signal array_obj_ref_728_index_offset_ack_1 : boolean;
  signal array_obj_ref_728_load_0_req_0 : boolean;
  signal array_obj_ref_728_load_0_ack_0 : boolean;
  signal array_obj_ref_728_load_0_req_1 : boolean;
  signal array_obj_ref_728_load_0_ack_1 : boolean;
  signal array_obj_ref_731_load_0_req_0 : boolean;
  signal array_obj_ref_731_load_0_ack_0 : boolean;
  signal array_obj_ref_731_load_0_req_1 : boolean;
  signal array_obj_ref_731_load_0_ack_1 : boolean;
  signal type_cast_733_inst_req_0 : boolean;
  signal type_cast_733_inst_ack_0 : boolean;
  signal type_cast_733_inst_req_1 : boolean;
  signal type_cast_733_inst_ack_1 : boolean;
  signal array_obj_ref_738_index_offset_req_0 : boolean;
  signal array_obj_ref_738_index_offset_ack_0 : boolean;
  signal array_obj_ref_738_index_offset_req_1 : boolean;
  signal array_obj_ref_738_index_offset_ack_1 : boolean;
  signal array_obj_ref_738_load_0_req_0 : boolean;
  signal array_obj_ref_738_load_0_ack_0 : boolean;
  signal array_obj_ref_738_load_0_req_1 : boolean;
  signal array_obj_ref_738_load_0_ack_1 : boolean;
  signal array_obj_ref_741_load_0_req_0 : boolean;
  signal array_obj_ref_741_load_0_ack_0 : boolean;
  signal array_obj_ref_741_load_0_req_1 : boolean;
  signal array_obj_ref_741_load_0_ack_1 : boolean;
  signal type_cast_743_inst_req_0 : boolean;
  signal type_cast_743_inst_ack_0 : boolean;
  signal type_cast_743_inst_req_1 : boolean;
  signal type_cast_743_inst_ack_1 : boolean;
  signal array_obj_ref_801_load_0_ack_0 : boolean;
  signal array_obj_ref_801_load_0_req_0 : boolean;
  signal array_obj_ref_748_index_offset_req_0 : boolean;
  signal array_obj_ref_748_index_offset_ack_0 : boolean;
  signal array_obj_ref_748_index_offset_req_1 : boolean;
  signal array_obj_ref_748_index_offset_ack_1 : boolean;
  signal array_obj_ref_748_load_0_req_0 : boolean;
  signal array_obj_ref_748_load_0_ack_0 : boolean;
  signal array_obj_ref_748_load_0_req_1 : boolean;
  signal array_obj_ref_748_load_0_ack_1 : boolean;
  signal array_obj_ref_751_load_0_req_0 : boolean;
  signal array_obj_ref_751_load_0_ack_0 : boolean;
  signal array_obj_ref_751_load_0_req_1 : boolean;
  signal array_obj_ref_751_load_0_ack_1 : boolean;
  signal type_cast_753_inst_req_0 : boolean;
  signal type_cast_753_inst_ack_0 : boolean;
  signal type_cast_753_inst_req_1 : boolean;
  signal type_cast_753_inst_ack_1 : boolean;
  signal array_obj_ref_758_index_offset_req_0 : boolean;
  signal array_obj_ref_758_index_offset_ack_0 : boolean;
  signal array_obj_ref_758_index_offset_req_1 : boolean;
  signal array_obj_ref_758_index_offset_ack_1 : boolean;
  signal array_obj_ref_758_load_0_req_0 : boolean;
  signal array_obj_ref_758_load_0_ack_0 : boolean;
  signal array_obj_ref_758_load_0_req_1 : boolean;
  signal array_obj_ref_758_load_0_ack_1 : boolean;
  signal array_obj_ref_761_load_0_req_0 : boolean;
  signal array_obj_ref_761_load_0_ack_0 : boolean;
  signal array_obj_ref_761_load_0_req_1 : boolean;
  signal array_obj_ref_761_load_0_ack_1 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_req_0 : boolean;
  signal array_obj_ref_768_index_offset_ack_0 : boolean;
  signal array_obj_ref_768_index_offset_req_1 : boolean;
  signal array_obj_ref_768_index_offset_ack_1 : boolean;
  signal array_obj_ref_768_load_0_req_0 : boolean;
  signal array_obj_ref_768_load_0_ack_0 : boolean;
  signal array_obj_ref_768_load_0_req_1 : boolean;
  signal array_obj_ref_768_load_0_ack_1 : boolean;
  signal array_obj_ref_771_load_0_req_0 : boolean;
  signal array_obj_ref_771_load_0_ack_0 : boolean;
  signal array_obj_ref_771_load_0_req_1 : boolean;
  signal array_obj_ref_771_load_0_ack_1 : boolean;
  signal type_cast_773_inst_req_0 : boolean;
  signal type_cast_773_inst_ack_0 : boolean;
  signal type_cast_773_inst_req_1 : boolean;
  signal type_cast_773_inst_ack_1 : boolean;
  signal array_obj_ref_778_index_offset_req_0 : boolean;
  signal array_obj_ref_778_index_offset_ack_0 : boolean;
  signal array_obj_ref_778_index_offset_req_1 : boolean;
  signal array_obj_ref_778_index_offset_ack_1 : boolean;
  signal array_obj_ref_778_load_0_req_0 : boolean;
  signal array_obj_ref_778_load_0_ack_0 : boolean;
  signal array_obj_ref_778_load_0_req_1 : boolean;
  signal array_obj_ref_778_load_0_ack_1 : boolean;
  signal array_obj_ref_781_load_0_req_0 : boolean;
  signal array_obj_ref_781_load_0_ack_0 : boolean;
  signal array_obj_ref_781_load_0_req_1 : boolean;
  signal array_obj_ref_781_load_0_ack_1 : boolean;
  signal type_cast_783_inst_req_0 : boolean;
  signal type_cast_783_inst_ack_0 : boolean;
  signal type_cast_783_inst_req_1 : boolean;
  signal type_cast_783_inst_ack_1 : boolean;
  signal array_obj_ref_788_index_offset_req_0 : boolean;
  signal array_obj_ref_788_index_offset_ack_0 : boolean;
  signal array_obj_ref_788_index_offset_req_1 : boolean;
  signal array_obj_ref_788_index_offset_ack_1 : boolean;
  signal array_obj_ref_788_load_0_req_0 : boolean;
  signal array_obj_ref_788_load_0_ack_0 : boolean;
  signal array_obj_ref_788_load_0_req_1 : boolean;
  signal array_obj_ref_788_load_0_ack_1 : boolean;
  signal array_obj_ref_791_load_0_req_0 : boolean;
  signal array_obj_ref_791_load_0_ack_0 : boolean;
  signal array_obj_ref_791_load_0_req_1 : boolean;
  signal array_obj_ref_791_load_0_ack_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal array_obj_ref_798_index_offset_req_0 : boolean;
  signal array_obj_ref_798_index_offset_ack_0 : boolean;
  signal array_obj_ref_798_index_offset_req_1 : boolean;
  signal array_obj_ref_798_index_offset_ack_1 : boolean;
  signal array_obj_ref_798_load_0_req_0 : boolean;
  signal array_obj_ref_798_load_0_ack_0 : boolean;
  signal array_obj_ref_808_index_offset_req_0 : boolean;
  signal array_obj_ref_808_index_offset_ack_0 : boolean;
  signal array_obj_ref_808_index_offset_req_1 : boolean;
  signal array_obj_ref_808_index_offset_ack_1 : boolean;
  signal array_obj_ref_808_load_0_req_0 : boolean;
  signal array_obj_ref_808_load_0_ack_0 : boolean;
  signal array_obj_ref_808_load_0_req_1 : boolean;
  signal array_obj_ref_808_load_0_ack_1 : boolean;
  signal array_obj_ref_811_load_0_req_0 : boolean;
  signal array_obj_ref_811_load_0_ack_0 : boolean;
  signal array_obj_ref_811_load_0_req_1 : boolean;
  signal array_obj_ref_811_load_0_ack_1 : boolean;
  signal type_cast_813_inst_req_0 : boolean;
  signal type_cast_813_inst_ack_0 : boolean;
  signal type_cast_813_inst_req_1 : boolean;
  signal type_cast_813_inst_ack_1 : boolean;
  signal array_obj_ref_818_index_offset_req_0 : boolean;
  signal array_obj_ref_818_index_offset_ack_0 : boolean;
  signal array_obj_ref_818_index_offset_req_1 : boolean;
  signal array_obj_ref_818_index_offset_ack_1 : boolean;
  signal array_obj_ref_818_load_0_req_0 : boolean;
  signal array_obj_ref_818_load_0_ack_0 : boolean;
  signal array_obj_ref_818_load_0_req_1 : boolean;
  signal array_obj_ref_818_load_0_ack_1 : boolean;
  signal array_obj_ref_821_load_0_req_0 : boolean;
  signal array_obj_ref_821_load_0_ack_0 : boolean;
  signal array_obj_ref_821_load_0_req_1 : boolean;
  signal array_obj_ref_821_load_0_ack_1 : boolean;
  signal type_cast_823_inst_req_0 : boolean;
  signal type_cast_823_inst_ack_0 : boolean;
  signal type_cast_823_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_1 : boolean;
  signal array_obj_ref_828_index_offset_req_0 : boolean;
  signal array_obj_ref_828_index_offset_ack_0 : boolean;
  signal array_obj_ref_828_index_offset_req_1 : boolean;
  signal array_obj_ref_828_index_offset_ack_1 : boolean;
  signal array_obj_ref_828_load_0_req_0 : boolean;
  signal array_obj_ref_828_load_0_ack_0 : boolean;
  signal array_obj_ref_828_load_0_req_1 : boolean;
  signal array_obj_ref_828_load_0_ack_1 : boolean;
  signal array_obj_ref_831_load_0_req_0 : boolean;
  signal array_obj_ref_831_load_0_ack_0 : boolean;
  signal array_obj_ref_831_load_0_req_1 : boolean;
  signal array_obj_ref_831_load_0_ack_1 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal type_cast_833_inst_req_1 : boolean;
  signal type_cast_833_inst_ack_1 : boolean;
  signal type_cast_839_inst_req_0 : boolean;
  signal type_cast_839_inst_ack_0 : boolean;
  signal type_cast_839_inst_req_1 : boolean;
  signal type_cast_839_inst_ack_1 : boolean;
  signal type_cast_845_inst_req_0 : boolean;
  signal type_cast_845_inst_ack_0 : boolean;
  signal type_cast_845_inst_req_1 : boolean;
  signal type_cast_845_inst_ack_1 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal type_cast_857_inst_req_0 : boolean;
  signal type_cast_857_inst_ack_0 : boolean;
  signal type_cast_857_inst_req_1 : boolean;
  signal type_cast_857_inst_ack_1 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_1 : boolean;
  signal type_cast_863_inst_ack_1 : boolean;
  signal type_cast_869_inst_req_0 : boolean;
  signal type_cast_869_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_1 : boolean;
  signal type_cast_869_inst_ack_1 : boolean;
  signal type_cast_875_inst_req_0 : boolean;
  signal type_cast_875_inst_ack_0 : boolean;
  signal type_cast_875_inst_req_1 : boolean;
  signal type_cast_875_inst_ack_1 : boolean;
  signal type_cast_881_inst_req_0 : boolean;
  signal type_cast_881_inst_ack_0 : boolean;
  signal type_cast_881_inst_req_1 : boolean;
  signal type_cast_881_inst_ack_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal type_cast_893_inst_req_0 : boolean;
  signal type_cast_893_inst_ack_0 : boolean;
  signal type_cast_893_inst_req_1 : boolean;
  signal type_cast_893_inst_ack_1 : boolean;
  signal type_cast_899_inst_req_0 : boolean;
  signal type_cast_899_inst_ack_0 : boolean;
  signal type_cast_899_inst_req_1 : boolean;
  signal type_cast_899_inst_ack_1 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal type_cast_911_inst_req_0 : boolean;
  signal type_cast_911_inst_ack_0 : boolean;
  signal type_cast_911_inst_req_1 : boolean;
  signal type_cast_911_inst_ack_1 : boolean;
  signal type_cast_917_inst_req_0 : boolean;
  signal type_cast_917_inst_ack_0 : boolean;
  signal type_cast_917_inst_req_1 : boolean;
  signal type_cast_917_inst_ack_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "mainAcc_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 13) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= I;
  I_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(10 downto 6) <= J;
  J_buffer <= in_buffer_data_out(10 downto 6);
  in_buffer_data_in(12 downto 11) <= col_to_be_replaced;
  col_to_be_replaced_buffer <= in_buffer_data_out(12 downto 11);
  in_buffer_data_in(tag_length + 12 downto 13) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 12 downto 13);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  mainAcc_CP_2438_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "mainAcc_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ofmap_pixel_buffer;
  ofmap_pixel <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mainAcc_CP_2438_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= mainAcc_CP_2438_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mainAcc_CP_2438_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,mainAcc_CP_2438_start,"mainAcc cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,mainAcc_CP_2438_symbol, "mainAcc cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  mainAcc_CP_2438: Block -- control-path 
    signal mainAcc_CP_2438_elements: BooleanArray(196 downto 0);
    -- 
  begin -- 
    mainAcc_CP_2438_elements(0) <= mainAcc_CP_2438_start;
    mainAcc_CP_2438_symbol <= mainAcc_CP_2438_elements(196);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	111 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	144 
    -- CP-element group 0: 	112 
    -- CP-element group 0: 	92 
    -- CP-element group 0: 	138 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	162 
    -- CP-element group 0: 	189 
    -- CP-element group 0: 	128 
    -- CP-element group 0: 	177 
    -- CP-element group 0: 	192 
    -- CP-element group 0: 	195 
    -- CP-element group 0: 	132 
    -- CP-element group 0: 	90 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	78 
    -- CP-element group 0: 	150 
    -- CP-element group 0: 	146 
    -- CP-element group 0: 	99 
    -- CP-element group 0: 	174 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	83 
    -- CP-element group 0: 	165 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	135 
    -- CP-element group 0: 	137 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	147 
    -- CP-element group 0: 	148 
    -- CP-element group 0: 	156 
    -- CP-element group 0: 	159 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	139 
    -- CP-element group 0: 	120 
    -- CP-element group 0: 	108 
    -- CP-element group 0: 	110 
    -- CP-element group 0: 	96 
    -- CP-element group 0: 	42 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	180 
    -- CP-element group 0: 	183 
    -- CP-element group 0: 	168 
    -- CP-element group 0: 	171 
    -- CP-element group 0: 	126 
    -- CP-element group 0: 	141 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	119 
    -- CP-element group 0: 	87 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	102 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	121 
    -- CP-element group 0: 	94 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	123 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	186 
    -- CP-element group 0: 	153 
    -- CP-element group 0: 	114 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	129 
    -- CP-element group 0: 	130 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	38 
    -- CP-element group 0:  members (485) 
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_computed_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_resized_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_resized_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_resized_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_computed_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_index_computed_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_root_address_calculated
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_start/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_complete/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_start/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_complete/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_start/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_complete/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_resized_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_computed_1
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_sample_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Update/cr
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_update_start_
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Update/$entry
      -- CP-element group 0: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Update/cr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_647_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_647_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_661_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_661_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_673_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_733_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_731_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_731_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_771_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_791_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_823_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_771_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_821_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_821_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_857_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_863_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_917_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_811_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_893_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_923_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_741_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_711_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_763_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_839_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_831_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_831_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_881_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_887_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_723_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_753_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_869_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_741_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_721_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_851_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_801_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_801_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_791_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_783_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_751_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_743_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_899_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_875_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_833_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_773_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_793_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_781_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_781_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_721_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_761_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_761_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_813_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_905_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_911_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_845_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_803_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_673_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_683_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_681_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_681_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_693_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_811_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_751_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_691_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_691_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_703_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_701_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_701_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_713_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_711_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_647_inst_req_1); -- 
    req_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_647_inst_req_0); -- 
    req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_661_inst_req_0); -- 
    req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_661_inst_req_1); -- 
    req_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_673_inst_req_0); -- 
    cr_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_733_inst_req_1); -- 
    cr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_718_load_0_req_1); -- 
    cr_3177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_731_load_0_req_1); -- 
    rr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_731_load_0_req_0); -- 
    rr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_771_load_0_req_0); -- 
    rr_3874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_791_load_0_req_0); -- 
    cr_4254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_823_inst_req_1); -- 
    cr_4205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_818_load_0_req_1); -- 
    cr_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_771_load_0_req_1); -- 
    req_4291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_828_index_offset_req_1); -- 
    req_3819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_788_index_offset_req_1); -- 
    cr_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_821_load_0_req_1); -- 
    rr_4228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_821_load_0_req_0); -- 
    req_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_758_index_offset_req_1); -- 
    cr_4428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_857_inst_req_1); -- 
    cr_4442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_863_inst_req_1); -- 
    cr_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_917_inst_req_1); -- 
    cr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_811_load_0_req_1); -- 
    cr_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_893_inst_req_1); -- 
    cr_4582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_923_inst_req_1); -- 
    req_3583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_768_index_offset_req_1); -- 
    req_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_798_index_offset_req_1); -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_741_load_0_req_1); -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_711_load_0_req_0); -- 
    req_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_728_index_offset_req_1); -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_778_index_offset_req_1); -- 
    cr_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_763_inst_req_1); -- 
    cr_4386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_839_inst_req_1); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_831_load_0_req_1); -- 
    rr_4346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_831_load_0_req_0); -- 
    cr_4484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_881_inst_req_1); -- 
    cr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_887_inst_req_1); -- 
    cr_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_723_inst_req_1); -- 
    cr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_753_inst_req_1); -- 
    cr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_748_load_0_req_1); -- 
    cr_4456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_869_inst_req_1); -- 
    rr_3284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_741_load_0_req_0); -- 
    rr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_721_load_0_req_0); -- 
    cr_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_778_load_0_req_1); -- 
    cr_4414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_851_inst_req_1); -- 
    cr_4003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_801_load_0_req_1); -- 
    rr_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_801_load_0_req_0); -- 
    cr_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_791_load_0_req_1); -- 
    cr_3782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_783_inst_req_1); -- 
    rr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_751_load_0_req_0); -- 
    req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_738_index_offset_req_1); -- 
    cr_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_743_inst_req_1); -- 
    cr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_738_load_0_req_1); -- 
    cr_3497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_758_load_0_req_1); -- 
    cr_4526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_899_inst_req_1); -- 
    cr_4470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_875_inst_req_1); -- 
    req_4055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_808_index_offset_req_1); -- 
    cr_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_833_inst_req_1); -- 
    cr_4323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_828_load_0_req_1); -- 
    req_2993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_718_index_offset_req_1); -- 
    cr_3664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_773_inst_req_1); -- 
    cr_3900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_793_inst_req_1); -- 
    cr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_788_load_0_req_1); -- 
    cr_3767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_781_load_0_req_1); -- 
    rr_3756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_781_load_0_req_0); -- 
    cr_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_721_load_0_req_1); -- 
    req_4173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_818_index_offset_req_1); -- 
    cr_3143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_728_load_0_req_1); -- 
    req_3347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_748_index_offset_req_1); -- 
    cr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_768_load_0_req_1); -- 
    cr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_761_load_0_req_1); -- 
    rr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_761_load_0_req_0); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_813_inst_req_1); -- 
    cr_4087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_808_load_0_req_1); -- 
    cr_4540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_905_inst_req_1); -- 
    cr_4554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_911_inst_req_1); -- 
    cr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_845_inst_req_1); -- 
    cr_4018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_803_inst_req_1); -- 
    cr_3969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_798_load_0_req_1); -- 
    req_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => MUX_673_inst_req_1); -- 
    cr_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_683_inst_req_1); -- 
    cr_2553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_678_load_0_req_1); -- 
    req_2516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_678_index_offset_req_0); -- 
    req_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_678_index_offset_req_1); -- 
    cr_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_681_load_0_req_1); -- 
    rr_2576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_681_load_0_req_0); -- 
    cr_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_693_inst_req_1); -- 
    cr_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_688_load_0_req_1); -- 
    rr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_811_load_0_req_0); -- 
    cr_3413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_751_load_0_req_1); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_688_index_offset_req_0); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_688_index_offset_req_1); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_691_load_0_req_1); -- 
    rr_2694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_691_load_0_req_0); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_703_inst_req_1); -- 
    cr_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_698_load_0_req_1); -- 
    req_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_698_index_offset_req_0); -- 
    req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_698_index_offset_req_1); -- 
    cr_2823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_701_load_0_req_1); -- 
    rr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_701_load_0_req_0); -- 
    cr_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => type_cast_713_inst_req_1); -- 
    cr_2907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_708_load_0_req_1); -- 
    req_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_708_index_offset_req_0); -- 
    req_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_708_index_offset_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(0), ack => array_obj_ref_711_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_sample_completed_
      -- CP-element group 1: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_start/$exit
      -- CP-element group 1: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_start/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_647_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_647_inst_ack_0, ack => mainAcc_CP_2438_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	44 
    -- CP-element group 2: 	53 
    -- CP-element group 2: 	62 
    -- CP-element group 2: 	71 
    -- CP-element group 2:  members (55) 
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_update_completed_
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_complete/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/MUX_647_complete/ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_resized_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_computed_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_resized_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_computed_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_resized_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_computed_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_resized_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_computed_1
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_647_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_647_inst_ack_1, ack => mainAcc_CP_2438_elements(2)); -- 
    req_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(2), ack => array_obj_ref_728_index_offset_req_0); -- 
    req_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(2), ack => array_obj_ref_718_index_offset_req_0); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(2), ack => array_obj_ref_748_index_offset_req_0); -- 
    req_3224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(2), ack => array_obj_ref_738_index_offset_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_sample_completed_
      -- CP-element group 3: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_start/$exit
      -- CP-element group 3: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_start/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_661_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_661_inst_ack_0, ack => mainAcc_CP_2438_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	80 
    -- CP-element group 4: 	89 
    -- CP-element group 4: 	98 
    -- CP-element group 4: 	107 
    -- CP-element group 4:  members (55) 
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_update_completed_
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_complete/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/MUX_661_complete/ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_resized_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_computed_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_resized_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_computed_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_resized_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_computed_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_resized_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_computed_1
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_661_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_661_inst_ack_1, ack => mainAcc_CP_2438_elements(4)); -- 
    req_3578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(4), ack => array_obj_ref_768_index_offset_req_0); -- 
    req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(4), ack => array_obj_ref_778_index_offset_req_0); -- 
    req_3814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(4), ack => array_obj_ref_788_index_offset_req_0); -- 
    req_3460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(4), ack => array_obj_ref_758_index_offset_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_sample_completed_
      -- CP-element group 5: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_start/$exit
      -- CP-element group 5: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_start/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_673_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_673_inst_ack_0, ack => mainAcc_CP_2438_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	143 
    -- CP-element group 6: 	116 
    -- CP-element group 6: 	125 
    -- CP-element group 6: 	134 
    -- CP-element group 6:  members (55) 
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_update_completed_
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_complete/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/MUX_673_complete/ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_resized_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_computed_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_resized_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_computed_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_resized_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_computed_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_resized_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_computed_1
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:MUX_673_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_673_inst_ack_1, ack => mainAcc_CP_2438_elements(6)); -- 
    req_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(6), ack => array_obj_ref_798_index_offset_req_0); -- 
    req_4050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(6), ack => array_obj_ref_808_index_offset_req_0); -- 
    req_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(6), ack => array_obj_ref_818_index_offset_req_0); -- 
    req_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(6), ack => array_obj_ref_828_index_offset_req_0); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	11 
    -- CP-element group 7: 	13 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	14 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_sample_start_
      -- CP-element group 7: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Sample/$entry
      -- CP-element group 7: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_683_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(7), ack => type_cast_683_inst_req_0); -- 
    mainAcc_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "mainAcc_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(11) & mainAcc_CP_2438_elements(13);
      gj_mainAcc_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	196 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_sample_complete
      -- CP-element group 8: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_offset_ack_0, ack => mainAcc_CP_2438_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (18) 
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_sample_start_
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_word_address_calculated
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_root_address_calculated
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_offset_calculated
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Update/$exit
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_final_index_sum_regn_Update/ack
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_base_plus_offset/$entry
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_base_plus_offset/$exit
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_base_plus_offset/sum_rename_req
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_base_plus_offset/sum_rename_ack
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_word_addrgen/$entry
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_word_addrgen/$exit
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_word_addrgen/root_register_req
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_word_addrgen/root_register_ack
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/$entry
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/word_0/$entry
      -- CP-element group 9: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_offset_ack_1, ack => mainAcc_CP_2438_elements(9)); -- 
    rr_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(9), ack => array_obj_ref_678_load_0_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_sample_completed_
      -- CP-element group 10: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/$exit
      -- CP-element group 10: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/$exit
      -- CP-element group 10: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_load_0_ack_0, ack => mainAcc_CP_2438_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	7 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_update_completed_
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/$exit
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/$exit
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/array_obj_ref_678_Merge/$entry
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/array_obj_ref_678_Merge/$exit
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/array_obj_ref_678_Merge/merge_req
      -- CP-element group 11: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_678_Update/array_obj_ref_678_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_678_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_load_0_ack_1, ack => mainAcc_CP_2438_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_sample_completed_
      -- CP-element group 12: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/$exit
      -- CP-element group 12: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_681_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_681_load_0_ack_0, ack => mainAcc_CP_2438_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	7 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_update_completed_
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/$exit
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/$exit
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/array_obj_ref_681_Merge/$entry
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/array_obj_ref_681_Merge/$exit
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/array_obj_ref_681_Merge/merge_req
      -- CP-element group 13: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_681_Update/array_obj_ref_681_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_681_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_681_load_0_ack_1, ack => mainAcc_CP_2438_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	7 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_sample_completed_
      -- CP-element group 14: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Sample/$exit
      -- CP-element group 14: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_683_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_0, ack => mainAcc_CP_2438_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	154 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_update_completed_
      -- CP-element group 15: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Update/$exit
      -- CP-element group 15: 	 assign_stmt_624_to_assign_stmt_924/type_cast_683_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_683_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_683_inst_ack_1, ack => mainAcc_CP_2438_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	22 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Sample/rr
      -- CP-element group 16: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_sample_start_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_693_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(16), ack => type_cast_693_inst_req_0); -- 
    mainAcc_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(20) & mainAcc_CP_2438_elements(22);
      gj_mainAcc_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	196 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Sample/ack
      -- CP-element group 17: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_0, ack => mainAcc_CP_2438_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (18) 
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/$entry
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/word_0/$entry
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_word_addrgen/$exit
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/word_0/rr
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_word_addrgen/root_register_ack
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_word_addrgen/root_register_req
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_word_addrgen/$entry
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_base_plus_offset/$exit
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_offset_calculated
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_base_plus_offset/$entry
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_sample_start_
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_word_address_calculated
      -- CP-element group 18: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_root_address_calculated
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_1, ack => mainAcc_CP_2438_elements(18)); -- 
    rr_2660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(18), ack => array_obj_ref_688_load_0_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/$exit
      -- CP-element group 19: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_sample_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_load_0_ack_0, ack => mainAcc_CP_2438_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/array_obj_ref_688_Merge/merge_ack
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/$exit
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/array_obj_ref_688_Merge/merge_req
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/$exit
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/array_obj_ref_688_Merge/$exit
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/array_obj_ref_688_Merge/$entry
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_688_update_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_688_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_load_0_ack_1, ack => mainAcc_CP_2438_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/word_0/ra
      -- CP-element group 21: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_sample_completed_
      -- CP-element group 21: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/$exit
      -- CP-element group 21: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_691_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_691_load_0_ack_0, ack => mainAcc_CP_2438_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	16 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/array_obj_ref_691_Merge/merge_req
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/array_obj_ref_691_Merge/$exit
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/array_obj_ref_691_Merge/$entry
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_update_completed_
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/array_obj_ref_691_Merge/merge_ack
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/word_access_complete/$exit
      -- CP-element group 22: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_691_Update/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_691_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_691_load_0_ack_1, ack => mainAcc_CP_2438_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Sample/ra
      -- CP-element group 23: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_sample_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_693_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_0, ack => mainAcc_CP_2438_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	160 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Update/$exit
      -- CP-element group 24: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_Update/ca
      -- CP-element group 24: 	 assign_stmt_624_to_assign_stmt_924/type_cast_693_update_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_693_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_1, ack => mainAcc_CP_2438_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	31 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Sample/rr
      -- CP-element group 25: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_sample_start_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_703_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(25), ack => type_cast_703_inst_req_0); -- 
    mainAcc_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(29) & mainAcc_CP_2438_elements(31);
      gj_mainAcc_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	196 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_sample_complete
      -- CP-element group 26: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Sample/$exit
      -- CP-element group 26: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_698_index_offset_ack_0, ack => mainAcc_CP_2438_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (18) 
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_root_address_calculated
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_word_addrgen/root_register_ack
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/$entry
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_word_address_calculated
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Update/$exit
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_offset_calculated
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_final_index_sum_regn_Update/ack
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_base_plus_offset/$entry
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_sample_start_
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/word_0/rr
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_base_plus_offset/$exit
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/word_0/$entry
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_word_addrgen/root_register_req
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_word_addrgen/$exit
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_word_addrgen/$entry
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_base_plus_offset/sum_rename_ack
      -- CP-element group 27: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_base_plus_offset/sum_rename_req
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_698_index_offset_ack_1, ack => mainAcc_CP_2438_elements(27)); -- 
    rr_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(27), ack => array_obj_ref_698_load_0_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_sample_completed_
      -- CP-element group 28: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/word_0/ra
      -- CP-element group 28: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/word_0/$exit
      -- CP-element group 28: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_698_load_0_ack_0, ack => mainAcc_CP_2438_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/array_obj_ref_698_Merge/$entry
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/array_obj_ref_698_Merge/$exit
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/array_obj_ref_698_Merge/merge_req
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/array_obj_ref_698_Merge/merge_ack
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/word_0/ca
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/$exit
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/$exit
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_update_completed_
      -- CP-element group 29: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_698_Update/word_access_complete/word_0/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_698_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_698_load_0_ack_1, ack => mainAcc_CP_2438_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/$exit
      -- CP-element group 30: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_sample_completed_
      -- CP-element group 30: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/$exit
      -- CP-element group 30: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/word_0/ra
      -- CP-element group 30: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_701_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_701_load_0_ack_0, ack => mainAcc_CP_2438_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	25 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/array_obj_ref_701_Merge/merge_ack
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/$exit
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/array_obj_ref_701_Merge/merge_req
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/array_obj_ref_701_Merge/$exit
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/$exit
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_update_completed_
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/word_access_complete/word_0/ca
      -- CP-element group 31: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_701_Update/array_obj_ref_701_Merge/$entry
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_701_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_701_load_0_ack_1, ack => mainAcc_CP_2438_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	25 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_sample_completed_
      -- CP-element group 32: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_703_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_0, ack => mainAcc_CP_2438_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	166 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_update_completed_
      -- CP-element group 33: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Update/$exit
      -- CP-element group 33: 	 assign_stmt_624_to_assign_stmt_924/type_cast_703_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_703_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_703_inst_ack_1, ack => mainAcc_CP_2438_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	38 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_sample_start_
      -- CP-element group 34: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_713_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(34), ack => type_cast_713_inst_req_0); -- 
    mainAcc_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(40) & mainAcc_CP_2438_elements(38);
      gj_mainAcc_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	196 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_sample_complete
      -- CP-element group 35: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_offset_ack_0, ack => mainAcc_CP_2438_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (18) 
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/word_0/rr
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_word_address_calculated
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_root_address_calculated
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_offset_calculated
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_base_plus_offset/sum_rename_req
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_base_plus_offset/$exit
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_base_plus_offset/sum_rename_ack
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Update/ack
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_word_addrgen/$entry
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_word_addrgen/$exit
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_word_addrgen/root_register_req
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_final_index_sum_regn_Update/$exit
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_word_addrgen/root_register_ack
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_sample_start_
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_base_plus_offset/$entry
      -- CP-element group 36: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/$entry
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_offset_ack_1, ack => mainAcc_CP_2438_elements(36)); -- 
    rr_2896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(36), ack => array_obj_ref_708_load_0_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_sample_completed_
      -- CP-element group 37: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/$exit
      -- CP-element group 37: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_load_0_ack_0, ack => mainAcc_CP_2438_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	34 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/array_obj_ref_708_Merge/$entry
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/$exit
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/array_obj_ref_708_Merge/$exit
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/array_obj_ref_708_Merge/merge_req
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/array_obj_ref_708_Merge/merge_ack
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_update_completed_
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/$exit
      -- CP-element group 38: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_708_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_708_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_load_0_ack_1, ack => mainAcc_CP_2438_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/$exit
      -- CP-element group 39: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_sample_completed_
      -- CP-element group 39: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/$exit
      -- CP-element group 39: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_711_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_711_load_0_ack_0, ack => mainAcc_CP_2438_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	34 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_update_completed_
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/word_0/$exit
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/$exit
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/array_obj_ref_711_Merge/merge_ack
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/array_obj_ref_711_Merge/merge_req
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/array_obj_ref_711_Merge/$exit
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/array_obj_ref_711_Merge/$entry
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/word_0/ca
      -- CP-element group 40: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_711_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_711_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_711_load_0_ack_1, ack => mainAcc_CP_2438_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_sample_completed_
      -- CP-element group 41: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Sample/$exit
      -- CP-element group 41: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_713_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_0, ack => mainAcc_CP_2438_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	0 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	172 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_update_completed_
      -- CP-element group 42: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Update/$exit
      -- CP-element group 42: 	 assign_stmt_624_to_assign_stmt_924/type_cast_713_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_713_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_713_inst_ack_1, ack => mainAcc_CP_2438_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	49 
    -- CP-element group 43: 	47 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	50 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_sample_start_
      -- CP-element group 43: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Sample/$entry
      -- CP-element group 43: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_723_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(43), ack => type_cast_723_inst_req_0); -- 
    mainAcc_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(49) & mainAcc_CP_2438_elements(47);
      gj_mainAcc_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	2 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	196 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_718_index_offset_ack_0, ack => mainAcc_CP_2438_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (18) 
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_sample_start_
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_word_address_calculated
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_root_address_calculated
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_offset_calculated
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_base_plus_offset/$entry
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_base_plus_offset/$exit
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_word_addrgen/$entry
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_word_addrgen/$exit
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_word_addrgen/root_register_req
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_word_addrgen/root_register_ack
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/$entry
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/$entry
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_718_index_offset_ack_1, ack => mainAcc_CP_2438_elements(45)); -- 
    rr_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(45), ack => array_obj_ref_718_load_0_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_sample_completed_
      -- CP-element group 46: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_718_load_0_ack_0, ack => mainAcc_CP_2438_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	43 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_update_completed_
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/$exit
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/array_obj_ref_718_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/array_obj_ref_718_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/array_obj_ref_718_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_718_Update/array_obj_ref_718_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_718_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_718_load_0_ack_1, ack => mainAcc_CP_2438_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_sample_completed_
      -- CP-element group 48: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/$exit
      -- CP-element group 48: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/$exit
      -- CP-element group 48: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_721_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_721_load_0_ack_0, ack => mainAcc_CP_2438_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	43 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_update_completed_
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/$exit
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/$exit
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/array_obj_ref_721_Merge/$entry
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/array_obj_ref_721_Merge/$exit
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/array_obj_ref_721_Merge/merge_req
      -- CP-element group 49: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_721_Update/array_obj_ref_721_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_721_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_721_load_0_ack_1, ack => mainAcc_CP_2438_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	43 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_sample_completed_
      -- CP-element group 50: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_723_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_723_inst_ack_0, ack => mainAcc_CP_2438_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	154 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_update_completed_
      -- CP-element group 51: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Update/$exit
      -- CP-element group 51: 	 assign_stmt_624_to_assign_stmt_924/type_cast_723_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_723_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_723_inst_ack_1, ack => mainAcc_CP_2438_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	58 
    -- CP-element group 52: 	56 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	59 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_sample_start_
      -- CP-element group 52: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_733_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(52), ack => type_cast_733_inst_req_0); -- 
    mainAcc_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(58) & mainAcc_CP_2438_elements(56);
      gj_mainAcc_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	2 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	196 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_sample_complete
      -- CP-element group 53: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Sample/$exit
      -- CP-element group 53: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_728_index_offset_ack_0, ack => mainAcc_CP_2438_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (18) 
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_sample_start_
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_word_address_calculated
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_root_address_calculated
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_offset_calculated
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Update/$exit
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_final_index_sum_regn_Update/ack
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_base_plus_offset/$entry
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_base_plus_offset/$exit
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_word_addrgen/$entry
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_word_addrgen/$exit
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_word_addrgen/root_register_req
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_word_addrgen/root_register_ack
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/$entry
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/$entry
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/word_0/$entry
      -- CP-element group 54: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_728_index_offset_ack_1, ack => mainAcc_CP_2438_elements(54)); -- 
    rr_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(54), ack => array_obj_ref_728_load_0_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_sample_completed_
      -- CP-element group 55: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/$exit
      -- CP-element group 55: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/$exit
      -- CP-element group 55: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/word_0/$exit
      -- CP-element group 55: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_728_load_0_ack_0, ack => mainAcc_CP_2438_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_update_completed_
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/$exit
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/$exit
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/word_0/$exit
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/word_access_complete/word_0/ca
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/array_obj_ref_728_Merge/$entry
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/array_obj_ref_728_Merge/$exit
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/array_obj_ref_728_Merge/merge_req
      -- CP-element group 56: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_728_Update/array_obj_ref_728_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_728_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_728_load_0_ack_1, ack => mainAcc_CP_2438_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_sample_completed_
      -- CP-element group 57: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/$exit
      -- CP-element group 57: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/$exit
      -- CP-element group 57: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/word_0/$exit
      -- CP-element group 57: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_731_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_731_load_0_ack_0, ack => mainAcc_CP_2438_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	52 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_update_completed_
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/$exit
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/$exit
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/word_0/$exit
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/word_access_complete/word_0/ca
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/array_obj_ref_731_Merge/$entry
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/array_obj_ref_731_Merge/$exit
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/array_obj_ref_731_Merge/merge_req
      -- CP-element group 58: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_731_Update/array_obj_ref_731_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_731_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_731_load_0_ack_1, ack => mainAcc_CP_2438_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	52 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_sample_completed_
      -- CP-element group 59: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Sample/$exit
      -- CP-element group 59: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_733_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_0, ack => mainAcc_CP_2438_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	160 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_update_completed_
      -- CP-element group 60: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Update/$exit
      -- CP-element group 60: 	 assign_stmt_624_to_assign_stmt_924/type_cast_733_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_733_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_1, ack => mainAcc_CP_2438_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	67 
    -- CP-element group 61: 	65 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	68 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_sample_start_
      -- CP-element group 61: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Sample/$entry
      -- CP-element group 61: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_743_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(61), ack => type_cast_743_inst_req_0); -- 
    mainAcc_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(67) & mainAcc_CP_2438_elements(65);
      gj_mainAcc_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	2 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	196 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_sample_complete
      -- CP-element group 62: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_index_offset_ack_0, ack => mainAcc_CP_2438_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/$entry
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_sample_start_
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_word_address_calculated
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_root_address_calculated
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_offset_calculated
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Update/$exit
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_final_index_sum_regn_Update/ack
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_base_plus_offset/$entry
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_base_plus_offset/$exit
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_word_addrgen/$entry
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_word_addrgen/$exit
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_word_addrgen/root_register_req
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_word_addrgen/root_register_ack
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/$entry
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_index_offset_ack_1, ack => mainAcc_CP_2438_elements(63)); -- 
    rr_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(63), ack => array_obj_ref_738_load_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_sample_completed_
      -- CP-element group 64: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/$exit
      -- CP-element group 64: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_load_0_ack_0, ack => mainAcc_CP_2438_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	61 
    -- CP-element group 65:  members (9) 
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_update_completed_
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/$exit
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/$exit
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/array_obj_ref_738_Merge/$entry
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/array_obj_ref_738_Merge/$exit
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/array_obj_ref_738_Merge/merge_req
      -- CP-element group 65: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_738_Update/array_obj_ref_738_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_738_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_load_0_ack_1, ack => mainAcc_CP_2438_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_sample_completed_
      -- CP-element group 66: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/$exit
      -- CP-element group 66: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/word_0/$exit
      -- CP-element group 66: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_741_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_741_load_0_ack_0, ack => mainAcc_CP_2438_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	61 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_update_completed_
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/$exit
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/$exit
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/word_0/$exit
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/word_access_complete/word_0/ca
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/array_obj_ref_741_Merge/$entry
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/array_obj_ref_741_Merge/$exit
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/array_obj_ref_741_Merge/merge_req
      -- CP-element group 67: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_741_Update/array_obj_ref_741_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_741_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_741_load_0_ack_1, ack => mainAcc_CP_2438_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	61 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_sample_completed_
      -- CP-element group 68: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Sample/$exit
      -- CP-element group 68: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_743_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_0, ack => mainAcc_CP_2438_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	166 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_update_completed_
      -- CP-element group 69: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Update/$exit
      -- CP-element group 69: 	 assign_stmt_624_to_assign_stmt_924/type_cast_743_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_743_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_1, ack => mainAcc_CP_2438_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	74 
    -- CP-element group 70: 	76 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	77 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_sample_start_
      -- CP-element group 70: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Sample/$entry
      -- CP-element group 70: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_753_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(70), ack => type_cast_753_inst_req_0); -- 
    mainAcc_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(74) & mainAcc_CP_2438_elements(76);
      gj_mainAcc_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	2 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	196 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_sample_complete
      -- CP-element group 71: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Sample/$exit
      -- CP-element group 71: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_index_offset_ack_0, ack => mainAcc_CP_2438_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (18) 
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_sample_start_
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_word_address_calculated
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_root_address_calculated
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_offset_calculated
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Update/$exit
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_final_index_sum_regn_Update/ack
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_base_plus_offset/$entry
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_base_plus_offset/$exit
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_word_addrgen/$entry
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_word_addrgen/$exit
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_word_addrgen/root_register_req
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_word_addrgen/root_register_ack
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/$entry
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_index_offset_ack_1, ack => mainAcc_CP_2438_elements(72)); -- 
    rr_3368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(72), ack => array_obj_ref_748_load_0_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_sample_completed_
      -- CP-element group 73: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/$exit
      -- CP-element group 73: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/$exit
      -- CP-element group 73: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/word_0/$exit
      -- CP-element group 73: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_load_0_ack_0, ack => mainAcc_CP_2438_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	70 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_update_completed_
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/$exit
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/$exit
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/word_0/$exit
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/word_access_complete/word_0/ca
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/array_obj_ref_748_Merge/$entry
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/array_obj_ref_748_Merge/$exit
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/array_obj_ref_748_Merge/merge_req
      -- CP-element group 74: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_748_Update/array_obj_ref_748_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_748_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_load_0_ack_1, ack => mainAcc_CP_2438_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_sample_completed_
      -- CP-element group 75: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/$exit
      -- CP-element group 75: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/$exit
      -- CP-element group 75: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/word_0/$exit
      -- CP-element group 75: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_751_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_751_load_0_ack_0, ack => mainAcc_CP_2438_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	70 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_update_completed_
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/$exit
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/$exit
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/word_0/$exit
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/word_access_complete/word_0/ca
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/array_obj_ref_751_Merge/$entry
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/array_obj_ref_751_Merge/$exit
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/array_obj_ref_751_Merge/merge_req
      -- CP-element group 76: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_751_Update/array_obj_ref_751_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_751_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_751_load_0_ack_1, ack => mainAcc_CP_2438_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	70 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_sample_completed_
      -- CP-element group 77: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Sample/$exit
      -- CP-element group 77: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_753_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_0, ack => mainAcc_CP_2438_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	0 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	172 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_update_completed_
      -- CP-element group 78: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Update/$exit
      -- CP-element group 78: 	 assign_stmt_624_to_assign_stmt_924/type_cast_753_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_753_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_1, ack => mainAcc_CP_2438_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	85 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_sample_start_
      -- CP-element group 79: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Sample/$entry
      -- CP-element group 79: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_763_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(79), ack => type_cast_763_inst_req_0); -- 
    mainAcc_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(83) & mainAcc_CP_2438_elements(85);
      gj_mainAcc_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	4 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	196 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_sample_complete
      -- CP-element group 80: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Sample/$exit
      -- CP-element group 80: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_index_offset_ack_0, ack => mainAcc_CP_2438_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (18) 
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_sample_start_
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_word_address_calculated
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_root_address_calculated
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_offset_calculated
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Update/$exit
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_final_index_sum_regn_Update/ack
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_base_plus_offset/$entry
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_base_plus_offset/$exit
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_base_plus_offset/sum_rename_req
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_base_plus_offset/sum_rename_ack
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_word_addrgen/$entry
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_word_addrgen/$exit
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_word_addrgen/root_register_req
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_word_addrgen/root_register_ack
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/$entry
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/$entry
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/word_0/$entry
      -- CP-element group 81: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_index_offset_ack_1, ack => mainAcc_CP_2438_elements(81)); -- 
    rr_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(81), ack => array_obj_ref_758_load_0_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_sample_completed_
      -- CP-element group 82: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/$exit
      -- CP-element group 82: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_load_0_ack_0, ack => mainAcc_CP_2438_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_update_completed_
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/$exit
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/$exit
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/array_obj_ref_758_Merge/$entry
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/array_obj_ref_758_Merge/$exit
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/array_obj_ref_758_Merge/merge_req
      -- CP-element group 83: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_758_Update/array_obj_ref_758_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_758_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_758_load_0_ack_1, ack => mainAcc_CP_2438_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_sample_completed_
      -- CP-element group 84: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/$exit
      -- CP-element group 84: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/$exit
      -- CP-element group 84: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_761_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_761_load_0_ack_0, ack => mainAcc_CP_2438_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	79 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_update_completed_
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/$exit
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/$exit
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/array_obj_ref_761_Merge/$entry
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/array_obj_ref_761_Merge/$exit
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/array_obj_ref_761_Merge/merge_req
      -- CP-element group 85: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_761_Update/array_obj_ref_761_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_761_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_761_load_0_ack_1, ack => mainAcc_CP_2438_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	79 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_sample_completed_
      -- CP-element group 86: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_763_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => mainAcc_CP_2438_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	0 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	151 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_update_completed_
      -- CP-element group 87: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Update/$exit
      -- CP-element group 87: 	 assign_stmt_624_to_assign_stmt_924/type_cast_763_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_763_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => mainAcc_CP_2438_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	92 
    -- CP-element group 88: 	94 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	95 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_sample_start_
      -- CP-element group 88: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_773_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(88), ack => type_cast_773_inst_req_0); -- 
    mainAcc_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(92) & mainAcc_CP_2438_elements(94);
      gj_mainAcc_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	4 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	196 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_sample_complete
      -- CP-element group 89: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Sample/$exit
      -- CP-element group 89: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_0, ack => mainAcc_CP_2438_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	0 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (18) 
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_sample_start_
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_word_address_calculated
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_root_address_calculated
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_offset_calculated
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Update/$exit
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_final_index_sum_regn_Update/ack
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_base_plus_offset/$entry
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_base_plus_offset/$exit
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_word_addrgen/$entry
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_word_addrgen/$exit
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_word_addrgen/root_register_req
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_word_addrgen/root_register_ack
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/$entry
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/$entry
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/word_0/$entry
      -- CP-element group 90: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_1, ack => mainAcc_CP_2438_elements(90)); -- 
    rr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(90), ack => array_obj_ref_768_load_0_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_sample_completed_
      -- CP-element group 91: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/$exit
      -- CP-element group 91: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_load_0_ack_0, ack => mainAcc_CP_2438_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	0 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	88 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_update_completed_
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/$exit
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/$exit
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/word_access_complete/word_0/ca
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/array_obj_ref_768_Merge/$entry
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/array_obj_ref_768_Merge/$exit
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/array_obj_ref_768_Merge/merge_req
      -- CP-element group 92: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_768_Update/array_obj_ref_768_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_768_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_load_0_ack_1, ack => mainAcc_CP_2438_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_sample_completed_
      -- CP-element group 93: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/$exit
      -- CP-element group 93: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_771_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_771_load_0_ack_0, ack => mainAcc_CP_2438_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	0 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	88 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_update_completed_
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/$exit
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/$exit
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/array_obj_ref_771_Merge/$entry
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/array_obj_ref_771_Merge/$exit
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/array_obj_ref_771_Merge/merge_req
      -- CP-element group 94: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_771_Update/array_obj_ref_771_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_771_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_771_load_0_ack_1, ack => mainAcc_CP_2438_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	88 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_sample_completed_
      -- CP-element group 95: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Sample/$exit
      -- CP-element group 95: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_773_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_773_inst_ack_0, ack => mainAcc_CP_2438_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	0 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	157 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_update_completed_
      -- CP-element group 96: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Update/$exit
      -- CP-element group 96: 	 assign_stmt_624_to_assign_stmt_924/type_cast_773_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_773_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_773_inst_ack_1, ack => mainAcc_CP_2438_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	101 
    -- CP-element group 97: 	103 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_sample_start_
      -- CP-element group 97: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Sample/$entry
      -- CP-element group 97: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_783_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(97), ack => type_cast_783_inst_req_0); -- 
    mainAcc_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(101) & mainAcc_CP_2438_elements(103);
      gj_mainAcc_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	4 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	196 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_sample_complete
      -- CP-element group 98: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_778_index_offset_ack_0, ack => mainAcc_CP_2438_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	0 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (18) 
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_sample_start_
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_word_address_calculated
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_root_address_calculated
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_offset_calculated
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Update/$exit
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_final_index_sum_regn_Update/ack
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_base_plus_offset/$entry
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_base_plus_offset/$exit
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_base_plus_offset/sum_rename_req
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_base_plus_offset/sum_rename_ack
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_word_addrgen/$entry
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_word_addrgen/$exit
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_word_addrgen/root_register_req
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_word_addrgen/root_register_ack
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/$entry
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/$entry
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/word_0/$entry
      -- CP-element group 99: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_778_index_offset_ack_1, ack => mainAcc_CP_2438_elements(99)); -- 
    rr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(99), ack => array_obj_ref_778_load_0_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_sample_completed_
      -- CP-element group 100: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/$exit
      -- CP-element group 100: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/$exit
      -- CP-element group 100: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/word_0/$exit
      -- CP-element group 100: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_778_load_0_ack_0, ack => mainAcc_CP_2438_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	97 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_update_completed_
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/$exit
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/$exit
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/word_0/$exit
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/word_access_complete/word_0/ca
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/array_obj_ref_778_Merge/$entry
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/array_obj_ref_778_Merge/$exit
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/array_obj_ref_778_Merge/merge_req
      -- CP-element group 101: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_778_Update/array_obj_ref_778_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_778_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_778_load_0_ack_1, ack => mainAcc_CP_2438_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	0 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_sample_completed_
      -- CP-element group 102: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/$exit
      -- CP-element group 102: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_781_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_load_0_ack_0, ack => mainAcc_CP_2438_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	97 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_update_completed_
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/$exit
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/$exit
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/array_obj_ref_781_Merge/$entry
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/array_obj_ref_781_Merge/$exit
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/array_obj_ref_781_Merge/merge_req
      -- CP-element group 103: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_781_Update/array_obj_ref_781_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_781_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_load_0_ack_1, ack => mainAcc_CP_2438_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_sample_completed_
      -- CP-element group 104: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Sample/$exit
      -- CP-element group 104: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_783_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_0, ack => mainAcc_CP_2438_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	163 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_update_completed_
      -- CP-element group 105: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Update/$exit
      -- CP-element group 105: 	 assign_stmt_624_to_assign_stmt_924/type_cast_783_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_783_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_1, ack => mainAcc_CP_2438_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	112 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	113 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_sample_start_
      -- CP-element group 106: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Sample/$entry
      -- CP-element group 106: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_793_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(106), ack => type_cast_793_inst_req_0); -- 
    mainAcc_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(112) & mainAcc_CP_2438_elements(110);
      gj_mainAcc_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	4 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	196 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_sample_complete
      -- CP-element group 107: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Sample/$exit
      -- CP-element group 107: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_788_index_offset_ack_0, ack => mainAcc_CP_2438_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	0 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (18) 
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_sample_start_
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_word_address_calculated
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_root_address_calculated
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_offset_calculated
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Update/$exit
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_final_index_sum_regn_Update/ack
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_base_plus_offset/$entry
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_base_plus_offset/$exit
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_base_plus_offset/sum_rename_req
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_base_plus_offset/sum_rename_ack
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_word_addrgen/$entry
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_word_addrgen/$exit
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_word_addrgen/root_register_req
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_word_addrgen/root_register_ack
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/$entry
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_788_index_offset_ack_1, ack => mainAcc_CP_2438_elements(108)); -- 
    rr_3840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(108), ack => array_obj_ref_788_load_0_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_sample_completed_
      -- CP-element group 109: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/$exit
      -- CP-element group 109: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/$exit
      -- CP-element group 109: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_788_load_0_ack_0, ack => mainAcc_CP_2438_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	0 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_update_completed_
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/$exit
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/$exit
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/array_obj_ref_788_Merge/$entry
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/array_obj_ref_788_Merge/$exit
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/array_obj_ref_788_Merge/merge_req
      -- CP-element group 110: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_788_Update/array_obj_ref_788_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_788_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_788_load_0_ack_1, ack => mainAcc_CP_2438_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	0 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_sample_completed_
      -- CP-element group 111: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/$exit
      -- CP-element group 111: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/$exit
      -- CP-element group 111: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_791_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_791_load_0_ack_0, ack => mainAcc_CP_2438_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	0 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	106 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_update_completed_
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/$exit
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/$exit
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/array_obj_ref_791_Merge/$entry
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/array_obj_ref_791_Merge/$exit
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/array_obj_ref_791_Merge/merge_req
      -- CP-element group 112: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_791_Update/array_obj_ref_791_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_791_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_791_load_0_ack_1, ack => mainAcc_CP_2438_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	106 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_sample_completed_
      -- CP-element group 113: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Sample/$exit
      -- CP-element group 113: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_793_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => mainAcc_CP_2438_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	0 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	169 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_update_completed_
      -- CP-element group 114: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Update/$exit
      -- CP-element group 114: 	 assign_stmt_624_to_assign_stmt_924/type_cast_793_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_793_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => mainAcc_CP_2438_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	119 
    -- CP-element group 115: 	121 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Sample/$entry
      -- CP-element group 115: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Sample/rr
      -- CP-element group 115: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_sample_start_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_803_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(115), ack => type_cast_803_inst_req_0); -- 
    mainAcc_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(119) & mainAcc_CP_2438_elements(121);
      gj_mainAcc_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	6 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	196 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_sample_complete
      -- CP-element group 116: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Sample/$exit
      -- CP-element group 116: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_index_offset_ack_0, ack => mainAcc_CP_2438_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (18) 
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_sample_start_
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_word_address_calculated
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_root_address_calculated
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_offset_calculated
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Update/$exit
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_final_index_sum_regn_Update/ack
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_base_plus_offset/$entry
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_base_plus_offset/$exit
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_base_plus_offset/sum_rename_req
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_base_plus_offset/sum_rename_ack
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_word_addrgen/$entry
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_word_addrgen/$exit
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_word_addrgen/root_register_req
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_word_addrgen/root_register_ack
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/$entry
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/$entry
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_index_offset_ack_1, ack => mainAcc_CP_2438_elements(117)); -- 
    rr_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(117), ack => array_obj_ref_798_load_0_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_sample_completed_
      -- CP-element group 118: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/$exit
      -- CP-element group 118: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/word_0/$exit
      -- CP-element group 118: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_load_0_ack_0, ack => mainAcc_CP_2438_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	0 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	115 
    -- CP-element group 119:  members (9) 
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/word_0/$exit
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/array_obj_ref_798_Merge/merge_ack
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/word_0/ca
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/array_obj_ref_798_Merge/merge_req
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/array_obj_ref_798_Merge/$entry
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/array_obj_ref_798_Merge/$exit
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/word_access_complete/$exit
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_update_completed_
      -- CP-element group 119: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_798_Update/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_798_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_load_0_ack_1, ack => mainAcc_CP_2438_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	0 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/$exit
      -- CP-element group 120: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_sample_completed_
      -- CP-element group 120: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/word_0/ra
      -- CP-element group 120: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_801_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_801_load_0_ack_0, ack => mainAcc_CP_2438_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	0 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	115 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/array_obj_ref_801_Merge/merge_ack
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/array_obj_ref_801_Merge/merge_req
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/array_obj_ref_801_Merge/$exit
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_update_completed_
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/array_obj_ref_801_Merge/$entry
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/word_access_complete/$exit
      -- CP-element group 121: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_801_Update/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_801_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_801_load_0_ack_1, ack => mainAcc_CP_2438_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Sample/ra
      -- CP-element group 122: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_sample_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_803_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_0, ack => mainAcc_CP_2438_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	0 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	151 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Update/ca
      -- CP-element group 123: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_Update/$exit
      -- CP-element group 123: 	 assign_stmt_624_to_assign_stmt_924/type_cast_803_update_completed_
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_803_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_1, ack => mainAcc_CP_2438_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	130 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_sample_start_
      -- CP-element group 124: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_813_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(124), ack => type_cast_813_inst_req_0); -- 
    mainAcc_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(128) & mainAcc_CP_2438_elements(130);
      gj_mainAcc_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	6 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	196 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_808_index_offset_ack_0, ack => mainAcc_CP_2438_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	0 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (18) 
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_word_address_calculated
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_sample_start_
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_root_address_calculated
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_offset_calculated
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_base_plus_offset/$entry
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_base_plus_offset/$exit
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_word_addrgen/$entry
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_word_addrgen/$exit
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_word_addrgen/root_register_req
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_word_addrgen/root_register_ack
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/$entry
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/$entry
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_808_index_offset_ack_1, ack => mainAcc_CP_2438_elements(126)); -- 
    rr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(126), ack => array_obj_ref_808_load_0_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_sample_completed_
      -- CP-element group 127: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/$exit
      -- CP-element group 127: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/$exit
      -- CP-element group 127: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/word_0/$exit
      -- CP-element group 127: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_808_load_0_ack_0, ack => mainAcc_CP_2438_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	0 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	124 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_update_completed_
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/$exit
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/$exit
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/word_0/$exit
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/word_access_complete/word_0/ca
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/array_obj_ref_808_Merge/$entry
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/array_obj_ref_808_Merge/$exit
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/array_obj_ref_808_Merge/merge_req
      -- CP-element group 128: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_808_Update/array_obj_ref_808_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_808_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_808_load_0_ack_1, ack => mainAcc_CP_2438_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	0 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_sample_completed_
      -- CP-element group 129: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/$exit
      -- CP-element group 129: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/$exit
      -- CP-element group 129: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/word_0/$exit
      -- CP-element group 129: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_811_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_811_load_0_ack_0, ack => mainAcc_CP_2438_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	0 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	124 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_update_completed_
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/$exit
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/$exit
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/word_0/$exit
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/word_access_complete/word_0/ca
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/array_obj_ref_811_Merge/$entry
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/array_obj_ref_811_Merge/$exit
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/array_obj_ref_811_Merge/merge_req
      -- CP-element group 130: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_811_Update/array_obj_ref_811_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_811_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_811_load_0_ack_1, ack => mainAcc_CP_2438_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	124 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_sample_completed_
      -- CP-element group 131: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Sample/$exit
      -- CP-element group 131: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_813_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_0, ack => mainAcc_CP_2438_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	0 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	157 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_update_completed_
      -- CP-element group 132: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Update/$exit
      -- CP-element group 132: 	 assign_stmt_624_to_assign_stmt_924/type_cast_813_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_813_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_1, ack => mainAcc_CP_2438_elements(132)); -- 
    -- CP-element group 133:  join  transition  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: 	139 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	140 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_sample_start_
      -- CP-element group 133: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Sample/$entry
      -- CP-element group 133: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_823_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(133), ack => type_cast_823_inst_req_0); -- 
    mainAcc_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(137) & mainAcc_CP_2438_elements(139);
      gj_mainAcc_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	6 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	196 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_sample_complete
      -- CP-element group 134: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_818_index_offset_ack_0, ack => mainAcc_CP_2438_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	0 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (18) 
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_sample_start_
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_word_address_calculated
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_root_address_calculated
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_offset_calculated
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Update/$exit
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_final_index_sum_regn_Update/ack
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_base_plus_offset/$entry
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_base_plus_offset/$exit
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_base_plus_offset/sum_rename_req
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_base_plus_offset/sum_rename_ack
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_word_addrgen/$entry
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_word_addrgen/$exit
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_word_addrgen/root_register_req
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_word_addrgen/root_register_ack
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/$entry
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/$entry
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/word_0/$entry
      -- CP-element group 135: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_818_index_offset_ack_1, ack => mainAcc_CP_2438_elements(135)); -- 
    rr_4194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(135), ack => array_obj_ref_818_load_0_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_sample_completed_
      -- CP-element group 136: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/$exit
      -- CP-element group 136: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/$exit
      -- CP-element group 136: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/word_0/$exit
      -- CP-element group 136: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_818_load_0_ack_0, ack => mainAcc_CP_2438_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	0 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (9) 
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_update_completed_
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/$exit
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/$exit
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/word_0/$exit
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/word_access_complete/word_0/ca
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/array_obj_ref_818_Merge/$entry
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/array_obj_ref_818_Merge/$exit
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/array_obj_ref_818_Merge/merge_req
      -- CP-element group 137: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_818_Update/array_obj_ref_818_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_818_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_818_load_0_ack_1, ack => mainAcc_CP_2438_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	0 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (5) 
      -- CP-element group 138: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_sample_completed_
      -- CP-element group 138: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/$exit
      -- CP-element group 138: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/word_0/$exit
      -- CP-element group 138: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_821_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_821_load_0_ack_0, ack => mainAcc_CP_2438_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	0 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	133 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_update_completed_
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/$exit
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/$exit
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/word_0/$exit
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/word_access_complete/word_0/ca
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/array_obj_ref_821_Merge/$entry
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/array_obj_ref_821_Merge/$exit
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/array_obj_ref_821_Merge/merge_req
      -- CP-element group 139: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_821_Update/array_obj_ref_821_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_821_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_821_load_0_ack_1, ack => mainAcc_CP_2438_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	133 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_sample_completed_
      -- CP-element group 140: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Sample/$exit
      -- CP-element group 140: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_823_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_0, ack => mainAcc_CP_2438_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	0 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	163 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_update_completed_
      -- CP-element group 141: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Update/$exit
      -- CP-element group 141: 	 assign_stmt_624_to_assign_stmt_924/type_cast_823_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_823_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_1, ack => mainAcc_CP_2438_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	146 
    -- CP-element group 142: 	148 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	149 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_sample_start_
      -- CP-element group 142: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Sample/$entry
      -- CP-element group 142: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_833_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(142), ack => type_cast_833_inst_req_0); -- 
    mainAcc_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(146) & mainAcc_CP_2438_elements(148);
      gj_mainAcc_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	6 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	196 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_sample_complete
      -- CP-element group 143: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Sample/$exit
      -- CP-element group 143: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_828_index_offset_ack_0, ack => mainAcc_CP_2438_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	0 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (18) 
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_sample_start_
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_word_address_calculated
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_root_address_calculated
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_offset_calculated
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Update/$exit
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_final_index_sum_regn_Update/ack
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_base_plus_offset/$entry
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_base_plus_offset/$exit
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_base_plus_offset/sum_rename_req
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_base_plus_offset/sum_rename_ack
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_word_addrgen/$entry
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_word_addrgen/$exit
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_word_addrgen/root_register_req
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_word_addrgen/root_register_ack
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/$entry
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/$entry
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/word_0/$entry
      -- CP-element group 144: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_828_index_offset_ack_1, ack => mainAcc_CP_2438_elements(144)); -- 
    rr_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(144), ack => array_obj_ref_828_load_0_req_0); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_sample_completed_
      -- CP-element group 145: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/$exit
      -- CP-element group 145: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/$exit
      -- CP-element group 145: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_828_load_0_ack_0, ack => mainAcc_CP_2438_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	0 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	142 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_update_completed_
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/$exit
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/$exit
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/array_obj_ref_828_Merge/$entry
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/array_obj_ref_828_Merge/$exit
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/array_obj_ref_828_Merge/merge_req
      -- CP-element group 146: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_828_Update/array_obj_ref_828_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_828_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_828_load_0_ack_1, ack => mainAcc_CP_2438_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	0 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_sample_completed_
      -- CP-element group 147: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/$exit
      -- CP-element group 147: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/$exit
      -- CP-element group 147: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/word_0/$exit
      -- CP-element group 147: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_831_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_831_load_0_ack_0, ack => mainAcc_CP_2438_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	0 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	142 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_update_completed_
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/$exit
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/$exit
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/word_0/$exit
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/word_access_complete/word_0/ca
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/array_obj_ref_831_Merge/$entry
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/array_obj_ref_831_Merge/$exit
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/array_obj_ref_831_Merge/merge_req
      -- CP-element group 148: 	 assign_stmt_624_to_assign_stmt_924/array_obj_ref_831_Update/array_obj_ref_831_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:array_obj_ref_831_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_831_load_0_ack_1, ack => mainAcc_CP_2438_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	142 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_sample_completed_
      -- CP-element group 149: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Sample/$exit
      -- CP-element group 149: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_833_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => mainAcc_CP_2438_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	0 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	169 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_update_completed_
      -- CP-element group 150: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Update/$exit
      -- CP-element group 150: 	 assign_stmt_624_to_assign_stmt_924/type_cast_833_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_833_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_1, ack => mainAcc_CP_2438_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	87 
    -- CP-element group 151: 	123 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_sample_start_
      -- CP-element group 151: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Sample/$entry
      -- CP-element group 151: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_839_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(151), ack => type_cast_839_inst_req_0); -- 
    mainAcc_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(87) & mainAcc_CP_2438_elements(123);
      gj_mainAcc_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_sample_completed_
      -- CP-element group 152: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Sample/$exit
      -- CP-element group 152: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_839_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_0, ack => mainAcc_CP_2438_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	0 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	175 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_update_completed_
      -- CP-element group 153: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Update/$exit
      -- CP-element group 153: 	 assign_stmt_624_to_assign_stmt_924/type_cast_839_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_839_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_1, ack => mainAcc_CP_2438_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	51 
    -- CP-element group 154: 	15 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_sample_start_
      -- CP-element group 154: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Sample/$entry
      -- CP-element group 154: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_845_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(154), ack => type_cast_845_inst_req_0); -- 
    mainAcc_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(51) & mainAcc_CP_2438_elements(15);
      gj_mainAcc_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_sample_completed_
      -- CP-element group 155: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Sample/$exit
      -- CP-element group 155: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_845_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_845_inst_ack_0, ack => mainAcc_CP_2438_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	0 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	175 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_update_completed_
      -- CP-element group 156: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Update/$exit
      -- CP-element group 156: 	 assign_stmt_624_to_assign_stmt_924/type_cast_845_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_845_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_845_inst_ack_1, ack => mainAcc_CP_2438_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	132 
    -- CP-element group 157: 	96 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_sample_start_
      -- CP-element group 157: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Sample/$entry
      -- CP-element group 157: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_851_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(157), ack => type_cast_851_inst_req_0); -- 
    mainAcc_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(132) & mainAcc_CP_2438_elements(96);
      gj_mainAcc_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_sample_completed_
      -- CP-element group 158: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Sample/$exit
      -- CP-element group 158: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_851_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => mainAcc_CP_2438_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	0 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	178 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_update_completed_
      -- CP-element group 159: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Update/$exit
      -- CP-element group 159: 	 assign_stmt_624_to_assign_stmt_924/type_cast_851_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_851_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => mainAcc_CP_2438_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	60 
    -- CP-element group 160: 	24 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_sample_start_
      -- CP-element group 160: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_857_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(160), ack => type_cast_857_inst_req_0); -- 
    mainAcc_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(60) & mainAcc_CP_2438_elements(24);
      gj_mainAcc_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_sample_completed_
      -- CP-element group 161: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Sample/$exit
      -- CP-element group 161: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_857_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_0, ack => mainAcc_CP_2438_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	0 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	178 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_update_completed_
      -- CP-element group 162: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Update/$exit
      -- CP-element group 162: 	 assign_stmt_624_to_assign_stmt_924/type_cast_857_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_857_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_1, ack => mainAcc_CP_2438_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	105 
    -- CP-element group 163: 	141 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_sample_start_
      -- CP-element group 163: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Sample/$entry
      -- CP-element group 163: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_863_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(163), ack => type_cast_863_inst_req_0); -- 
    mainAcc_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(105) & mainAcc_CP_2438_elements(141);
      gj_mainAcc_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_sample_completed_
      -- CP-element group 164: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Sample/$exit
      -- CP-element group 164: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_863_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => mainAcc_CP_2438_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	0 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	181 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_update_completed_
      -- CP-element group 165: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Update/$exit
      -- CP-element group 165: 	 assign_stmt_624_to_assign_stmt_924/type_cast_863_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_863_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_1, ack => mainAcc_CP_2438_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	69 
    -- CP-element group 166: 	33 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_sample_start_
      -- CP-element group 166: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Sample/$entry
      -- CP-element group 166: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_869_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(166), ack => type_cast_869_inst_req_0); -- 
    mainAcc_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(69) & mainAcc_CP_2438_elements(33);
      gj_mainAcc_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_sample_completed_
      -- CP-element group 167: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Sample/$exit
      -- CP-element group 167: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_869_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_0, ack => mainAcc_CP_2438_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	0 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	181 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_update_completed_
      -- CP-element group 168: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Update/$exit
      -- CP-element group 168: 	 assign_stmt_624_to_assign_stmt_924/type_cast_869_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_869_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_1, ack => mainAcc_CP_2438_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	150 
    -- CP-element group 169: 	114 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_sample_start_
      -- CP-element group 169: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Sample/$entry
      -- CP-element group 169: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_875_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(169), ack => type_cast_875_inst_req_0); -- 
    mainAcc_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(150) & mainAcc_CP_2438_elements(114);
      gj_mainAcc_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_sample_completed_
      -- CP-element group 170: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Sample/$exit
      -- CP-element group 170: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_875_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_875_inst_ack_0, ack => mainAcc_CP_2438_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	0 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	184 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_update_completed_
      -- CP-element group 171: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Update/$exit
      -- CP-element group 171: 	 assign_stmt_624_to_assign_stmt_924/type_cast_875_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_875_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_875_inst_ack_1, ack => mainAcc_CP_2438_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	78 
    -- CP-element group 172: 	42 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_sample_start_
      -- CP-element group 172: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_881_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(172), ack => type_cast_881_inst_req_0); -- 
    mainAcc_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(78) & mainAcc_CP_2438_elements(42);
      gj_mainAcc_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_sample_completed_
      -- CP-element group 173: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Sample/$exit
      -- CP-element group 173: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_881_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_881_inst_ack_0, ack => mainAcc_CP_2438_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	0 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	184 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_update_completed_
      -- CP-element group 174: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Update/$exit
      -- CP-element group 174: 	 assign_stmt_624_to_assign_stmt_924/type_cast_881_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_881_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_881_inst_ack_1, ack => mainAcc_CP_2438_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	156 
    -- CP-element group 175: 	153 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_sample_start_
      -- CP-element group 175: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Sample/$entry
      -- CP-element group 175: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_887_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(175), ack => type_cast_887_inst_req_0); -- 
    mainAcc_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(156) & mainAcc_CP_2438_elements(153);
      gj_mainAcc_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_sample_completed_
      -- CP-element group 176: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Sample/$exit
      -- CP-element group 176: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_887_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => mainAcc_CP_2438_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	0 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	187 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_update_completed_
      -- CP-element group 177: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Update/$exit
      -- CP-element group 177: 	 assign_stmt_624_to_assign_stmt_924/type_cast_887_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_887_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => mainAcc_CP_2438_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	162 
    -- CP-element group 178: 	159 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_sample_start_
      -- CP-element group 178: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Sample/$entry
      -- CP-element group 178: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_893_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(178), ack => type_cast_893_inst_req_0); -- 
    mainAcc_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(162) & mainAcc_CP_2438_elements(159);
      gj_mainAcc_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_sample_completed_
      -- CP-element group 179: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Sample/$exit
      -- CP-element group 179: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_893_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_0, ack => mainAcc_CP_2438_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	0 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	187 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_update_completed_
      -- CP-element group 180: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Update/$exit
      -- CP-element group 180: 	 assign_stmt_624_to_assign_stmt_924/type_cast_893_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_893_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_1, ack => mainAcc_CP_2438_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	165 
    -- CP-element group 181: 	168 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_sample_start_
      -- CP-element group 181: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Sample/$entry
      -- CP-element group 181: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_899_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(181), ack => type_cast_899_inst_req_0); -- 
    mainAcc_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(165) & mainAcc_CP_2438_elements(168);
      gj_mainAcc_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_sample_completed_
      -- CP-element group 182: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Sample/$exit
      -- CP-element group 182: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_899_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_0, ack => mainAcc_CP_2438_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	0 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	190 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_update_completed_
      -- CP-element group 183: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Update/$exit
      -- CP-element group 183: 	 assign_stmt_624_to_assign_stmt_924/type_cast_899_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_899_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_1, ack => mainAcc_CP_2438_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	174 
    -- CP-element group 184: 	171 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_sample_start_
      -- CP-element group 184: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Sample/$entry
      -- CP-element group 184: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_905_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(184), ack => type_cast_905_inst_req_0); -- 
    mainAcc_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(174) & mainAcc_CP_2438_elements(171);
      gj_mainAcc_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_sample_completed_
      -- CP-element group 185: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Sample/$exit
      -- CP-element group 185: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_905_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => mainAcc_CP_2438_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	0 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	190 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_update_completed_
      -- CP-element group 186: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Update/$exit
      -- CP-element group 186: 	 assign_stmt_624_to_assign_stmt_924/type_cast_905_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_905_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => mainAcc_CP_2438_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	177 
    -- CP-element group 187: 	180 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_sample_start_
      -- CP-element group 187: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Sample/$entry
      -- CP-element group 187: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_911_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(187), ack => type_cast_911_inst_req_0); -- 
    mainAcc_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(177) & mainAcc_CP_2438_elements(180);
      gj_mainAcc_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_sample_completed_
      -- CP-element group 188: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Sample/$exit
      -- CP-element group 188: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_911_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_911_inst_ack_0, ack => mainAcc_CP_2438_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	0 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	193 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_update_completed_
      -- CP-element group 189: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Update/$exit
      -- CP-element group 189: 	 assign_stmt_624_to_assign_stmt_924/type_cast_911_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_911_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_911_inst_ack_1, ack => mainAcc_CP_2438_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	183 
    -- CP-element group 190: 	186 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_sample_start_
      -- CP-element group 190: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Sample/$entry
      -- CP-element group 190: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_917_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(190), ack => type_cast_917_inst_req_0); -- 
    mainAcc_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(183) & mainAcc_CP_2438_elements(186);
      gj_mainAcc_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_sample_completed_
      -- CP-element group 191: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Sample/$exit
      -- CP-element group 191: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_917_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_917_inst_ack_0, ack => mainAcc_CP_2438_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	0 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_update_completed_
      -- CP-element group 192: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Update/$exit
      -- CP-element group 192: 	 assign_stmt_624_to_assign_stmt_924/type_cast_917_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_917_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_917_inst_ack_1, ack => mainAcc_CP_2438_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	189 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_sample_start_
      -- CP-element group 193: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Sample/$entry
      -- CP-element group 193: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Sample/rr
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_923_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc_CP_2438_elements(193), ack => type_cast_923_inst_req_0); -- 
    mainAcc_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(189) & mainAcc_CP_2438_elements(192);
      gj_mainAcc_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_sample_completed_
      -- CP-element group 194: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Sample/ra
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_923_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => mainAcc_CP_2438_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	0 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_update_completed_
      -- CP-element group 195: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Update/$exit
      -- CP-element group 195: 	 assign_stmt_624_to_assign_stmt_924/type_cast_923_Update/ca
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:type_cast_923_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => mainAcc_CP_2438_elements(195)); -- 
    -- CP-element group 196:  join  transition  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	143 
    -- CP-element group 196: 	80 
    -- CP-element group 196: 	44 
    -- CP-element group 196: 	195 
    -- CP-element group 196: 	89 
    -- CP-element group 196: 	116 
    -- CP-element group 196: 	98 
    -- CP-element group 196: 	53 
    -- CP-element group 196: 	107 
    -- CP-element group 196: 	62 
    -- CP-element group 196: 	125 
    -- CP-element group 196: 	134 
    -- CP-element group 196: 	71 
    -- CP-element group 196: 	8 
    -- CP-element group 196: 	17 
    -- CP-element group 196: 	26 
    -- CP-element group 196: 	35 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 $exit
      -- CP-element group 196: 	 assign_stmt_624_to_assign_stmt_924/$exit
      -- 
    -- logger for CP element group mainAcc_CP_2438_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc_CP_2438_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc:CP:mainAcc_CP_2438_elements(196) fired."); 
        -- 
      end if; --
    end process; 
    mainAcc_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "mainAcc_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= mainAcc_CP_2438_elements(143) & mainAcc_CP_2438_elements(80) & mainAcc_CP_2438_elements(44) & mainAcc_CP_2438_elements(195) & mainAcc_CP_2438_elements(89) & mainAcc_CP_2438_elements(116) & mainAcc_CP_2438_elements(98) & mainAcc_CP_2438_elements(53) & mainAcc_CP_2438_elements(107) & mainAcc_CP_2438_elements(62) & mainAcc_CP_2438_elements(125) & mainAcc_CP_2438_elements(134) & mainAcc_CP_2438_elements(71) & mainAcc_CP_2438_elements(8) & mainAcc_CP_2438_elements(17) & mainAcc_CP_2438_elements(26) & mainAcc_CP_2438_elements(35);
      gj_mainAcc_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc_CP_2438_elements(196), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_838_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_844_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_850_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_856_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_862_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_868_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_874_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_880_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_886_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_892_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_898_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_904_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_910_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_916_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_922_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_659_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_671_wire : std_logic_vector(1 downto 0);
    signal EQ_u2_u1_640_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_666_wire : std_logic_vector(0 downto 0);
    signal MUL_u16_u16_682_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_692_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_702_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_712_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_722_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_732_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_742_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_752_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_762_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_772_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_782_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_792_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_802_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_812_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_822_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_832_wire : std_logic_vector(15 downto 0);
    signal R_col_to_be_replaced_1_717_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_717_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_727_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_727_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_737_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_737_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_747_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_747_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_757_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_757_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_767_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_767_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_777_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_777_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_787_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_787_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_797_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_797_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_807_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_807_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_817_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_817_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_827_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_827_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_677_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_677_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_687_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_687_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_697_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_697_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_707_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_707_scaled : std_logic_vector(3 downto 0);
    signal SUB_u2_u2_645_wire : std_logic_vector(1 downto 0);
    signal SUB_u2_u2_655_wire : std_logic_vector(1 downto 0);
    signal UGE_u2_u1_652_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_678_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_678_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_678_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_678_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_681_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_681_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_681_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_688_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_688_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_688_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_691_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_691_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_691_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_698_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_698_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_698_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_701_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_701_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_701_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_708_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_708_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_708_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_711_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_711_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_711_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_718_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_718_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_718_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_721_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_721_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_721_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_728_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_728_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_728_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_731_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_731_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_731_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_738_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_738_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_738_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_741_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_741_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_741_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_748_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_748_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_748_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_751_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_751_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_751_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_758_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_758_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_758_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_761_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_761_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_761_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_768_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_768_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_768_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_771_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_771_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_771_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_778_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_778_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_778_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_781_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_781_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_781_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_788_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_788_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_788_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_791_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_791_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_791_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_798_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_798_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_798_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_801_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_801_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_801_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_808_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_808_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_808_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_811_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_811_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_811_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_818_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_818_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_818_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_821_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_821_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_821_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_828_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_828_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_828_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_831_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_831_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_831_word_address_0 : std_logic_vector(3 downto 0);
    signal col_to_be_replaced_1_648 : std_logic_vector(1 downto 0);
    signal col_to_be_replaced_2_662 : std_logic_vector(1 downto 0);
    signal col_to_be_replaced_3_674 : std_logic_vector(1 downto 0);
    signal konst_639_wire_constant : std_logic_vector(1 downto 0);
    signal konst_644_wire_constant : std_logic_vector(1 downto 0);
    signal konst_651_wire_constant : std_logic_vector(1 downto 0);
    signal konst_654_wire_constant : std_logic_vector(1 downto 0);
    signal konst_658_wire_constant : std_logic_vector(1 downto 0);
    signal konst_665_wire_constant : std_logic_vector(1 downto 0);
    signal konst_670_wire_constant : std_logic_vector(1 downto 0);
    signal one_628 : std_logic_vector(1 downto 0);
    signal pp00_804 : std_logic_vector(15 downto 0);
    signal pp01_764 : std_logic_vector(15 downto 0);
    signal pp02_724 : std_logic_vector(15 downto 0);
    signal pp03_684 : std_logic_vector(15 downto 0);
    signal pp10_814 : std_logic_vector(15 downto 0);
    signal pp11_774 : std_logic_vector(15 downto 0);
    signal pp12_734 : std_logic_vector(15 downto 0);
    signal pp13_694 : std_logic_vector(15 downto 0);
    signal pp20_824 : std_logic_vector(15 downto 0);
    signal pp21_784 : std_logic_vector(15 downto 0);
    signal pp22_744 : std_logic_vector(15 downto 0);
    signal pp23_704 : std_logic_vector(15 downto 0);
    signal pp30_834 : std_logic_vector(15 downto 0);
    signal pp31_794 : std_logic_vector(15 downto 0);
    signal pp32_754 : std_logic_vector(15 downto 0);
    signal pp33_714 : std_logic_vector(15 downto 0);
    signal sum0_840 : std_logic_vector(15 downto 0);
    signal sum10_888 : std_logic_vector(15 downto 0);
    signal sum11_894 : std_logic_vector(15 downto 0);
    signal sum12_900 : std_logic_vector(15 downto 0);
    signal sum13_906 : std_logic_vector(15 downto 0);
    signal sum1_846 : std_logic_vector(15 downto 0);
    signal sum20_912 : std_logic_vector(15 downto 0);
    signal sum21_918 : std_logic_vector(15 downto 0);
    signal sum2_852 : std_logic_vector(15 downto 0);
    signal sum3_858 : std_logic_vector(15 downto 0);
    signal sum4_864 : std_logic_vector(15 downto 0);
    signal sum5_870 : std_logic_vector(15 downto 0);
    signal sum6_876 : std_logic_vector(15 downto 0);
    signal sum7_882 : std_logic_vector(15 downto 0);
    signal three_636 : std_logic_vector(1 downto 0);
    signal two_632 : std_logic_vector(1 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_646_wire : std_logic_vector(1 downto 0);
    signal type_cast_656_wire : std_logic_vector(1 downto 0);
    signal type_cast_660_wire : std_logic_vector(1 downto 0);
    signal type_cast_668_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_672_wire : std_logic_vector(1 downto 0);
    signal zero_624 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_678_constant_part_of_offset <= "0000";
    array_obj_ref_678_offset_scale_factor_0 <= "0100";
    array_obj_ref_678_offset_scale_factor_1 <= "0001";
    array_obj_ref_678_resized_base_address <= "0000";
    array_obj_ref_678_word_offset_0 <= "0000";
    array_obj_ref_681_word_address_0 <= "0011";
    array_obj_ref_688_constant_part_of_offset <= "0100";
    array_obj_ref_688_offset_scale_factor_0 <= "0100";
    array_obj_ref_688_offset_scale_factor_1 <= "0001";
    array_obj_ref_688_resized_base_address <= "0000";
    array_obj_ref_688_word_offset_0 <= "0000";
    array_obj_ref_691_word_address_0 <= "0111";
    array_obj_ref_698_constant_part_of_offset <= "1000";
    array_obj_ref_698_offset_scale_factor_0 <= "0100";
    array_obj_ref_698_offset_scale_factor_1 <= "0001";
    array_obj_ref_698_resized_base_address <= "0000";
    array_obj_ref_698_word_offset_0 <= "0000";
    array_obj_ref_701_word_address_0 <= "1011";
    array_obj_ref_708_constant_part_of_offset <= "1100";
    array_obj_ref_708_offset_scale_factor_0 <= "0100";
    array_obj_ref_708_offset_scale_factor_1 <= "0001";
    array_obj_ref_708_resized_base_address <= "0000";
    array_obj_ref_708_word_offset_0 <= "0000";
    array_obj_ref_711_word_address_0 <= "1111";
    array_obj_ref_718_constant_part_of_offset <= "0000";
    array_obj_ref_718_offset_scale_factor_0 <= "0100";
    array_obj_ref_718_offset_scale_factor_1 <= "0001";
    array_obj_ref_718_resized_base_address <= "0000";
    array_obj_ref_718_word_offset_0 <= "0000";
    array_obj_ref_721_word_address_0 <= "0010";
    array_obj_ref_728_constant_part_of_offset <= "0100";
    array_obj_ref_728_offset_scale_factor_0 <= "0100";
    array_obj_ref_728_offset_scale_factor_1 <= "0001";
    array_obj_ref_728_resized_base_address <= "0000";
    array_obj_ref_728_word_offset_0 <= "0000";
    array_obj_ref_731_word_address_0 <= "0110";
    array_obj_ref_738_constant_part_of_offset <= "1000";
    array_obj_ref_738_offset_scale_factor_0 <= "0100";
    array_obj_ref_738_offset_scale_factor_1 <= "0001";
    array_obj_ref_738_resized_base_address <= "0000";
    array_obj_ref_738_word_offset_0 <= "0000";
    array_obj_ref_741_word_address_0 <= "1010";
    array_obj_ref_748_constant_part_of_offset <= "1100";
    array_obj_ref_748_offset_scale_factor_0 <= "0100";
    array_obj_ref_748_offset_scale_factor_1 <= "0001";
    array_obj_ref_748_resized_base_address <= "0000";
    array_obj_ref_748_word_offset_0 <= "0000";
    array_obj_ref_751_word_address_0 <= "1110";
    array_obj_ref_758_constant_part_of_offset <= "0000";
    array_obj_ref_758_offset_scale_factor_0 <= "0100";
    array_obj_ref_758_offset_scale_factor_1 <= "0001";
    array_obj_ref_758_resized_base_address <= "0000";
    array_obj_ref_758_word_offset_0 <= "0000";
    array_obj_ref_761_word_address_0 <= "0001";
    array_obj_ref_768_constant_part_of_offset <= "0100";
    array_obj_ref_768_offset_scale_factor_0 <= "0100";
    array_obj_ref_768_offset_scale_factor_1 <= "0001";
    array_obj_ref_768_resized_base_address <= "0000";
    array_obj_ref_768_word_offset_0 <= "0000";
    array_obj_ref_771_word_address_0 <= "0101";
    array_obj_ref_778_constant_part_of_offset <= "1000";
    array_obj_ref_778_offset_scale_factor_0 <= "0100";
    array_obj_ref_778_offset_scale_factor_1 <= "0001";
    array_obj_ref_778_resized_base_address <= "0000";
    array_obj_ref_778_word_offset_0 <= "0000";
    array_obj_ref_781_word_address_0 <= "1001";
    array_obj_ref_788_constant_part_of_offset <= "1100";
    array_obj_ref_788_offset_scale_factor_0 <= "0100";
    array_obj_ref_788_offset_scale_factor_1 <= "0001";
    array_obj_ref_788_resized_base_address <= "0000";
    array_obj_ref_788_word_offset_0 <= "0000";
    array_obj_ref_791_word_address_0 <= "1101";
    array_obj_ref_798_constant_part_of_offset <= "0000";
    array_obj_ref_798_offset_scale_factor_0 <= "0100";
    array_obj_ref_798_offset_scale_factor_1 <= "0001";
    array_obj_ref_798_resized_base_address <= "0000";
    array_obj_ref_798_word_offset_0 <= "0000";
    array_obj_ref_801_word_address_0 <= "0000";
    array_obj_ref_808_constant_part_of_offset <= "0100";
    array_obj_ref_808_offset_scale_factor_0 <= "0100";
    array_obj_ref_808_offset_scale_factor_1 <= "0001";
    array_obj_ref_808_resized_base_address <= "0000";
    array_obj_ref_808_word_offset_0 <= "0000";
    array_obj_ref_811_word_address_0 <= "0100";
    array_obj_ref_818_constant_part_of_offset <= "1000";
    array_obj_ref_818_offset_scale_factor_0 <= "0100";
    array_obj_ref_818_offset_scale_factor_1 <= "0001";
    array_obj_ref_818_resized_base_address <= "0000";
    array_obj_ref_818_word_offset_0 <= "0000";
    array_obj_ref_821_word_address_0 <= "1000";
    array_obj_ref_828_constant_part_of_offset <= "1100";
    array_obj_ref_828_offset_scale_factor_0 <= "0100";
    array_obj_ref_828_offset_scale_factor_1 <= "0001";
    array_obj_ref_828_resized_base_address <= "0000";
    array_obj_ref_828_word_offset_0 <= "0000";
    array_obj_ref_831_word_address_0 <= "1100";
    konst_639_wire_constant <= "00";
    konst_644_wire_constant <= "01";
    konst_651_wire_constant <= "10";
    konst_654_wire_constant <= "10";
    konst_658_wire_constant <= "10";
    konst_665_wire_constant <= "11";
    konst_670_wire_constant <= "01";
    one_628 <= "01";
    three_636 <= "11";
    two_632 <= "10";
    type_cast_642_wire_constant <= "11";
    type_cast_668_wire_constant <= "00";
    zero_624 <= "00";
    -- logger for split-operator MUX_647_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_647_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_647_inst:started:   inputs: " & " EQ_u2_u1_640_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_640_wire) & " type_cast_642_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_642_wire_constant) & " type_cast_646_wire = "& Convert_SLV_To_Hex_String(type_cast_646_wire));
          --
        end if; 
        if MUX_647_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_647_inst:finished:  outputs: " & " col_to_be_replaced_1_648= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_1_648));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_647_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_647_inst_req_0;
      MUX_647_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_647_inst_req_1;
      MUX_647_inst_ack_1<= update_ack(0);
      MUX_647_inst: SelectSplitProtocol generic map(name => "MUX_647_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_642_wire_constant, y => type_cast_646_wire, sel => EQ_u2_u1_640_wire, z => col_to_be_replaced_1_648, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_661_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_661_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_661_inst:started:   inputs: " & " UGE_u2_u1_652_wire = "& Convert_SLV_To_Hex_String(UGE_u2_u1_652_wire) & " type_cast_656_wire = "& Convert_SLV_To_Hex_String(type_cast_656_wire) & " type_cast_660_wire = "& Convert_SLV_To_Hex_String(type_cast_660_wire));
          --
        end if; 
        if MUX_661_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_661_inst:finished:  outputs: " & " col_to_be_replaced_2_662= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_2_662));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_661_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_661_inst_req_0;
      MUX_661_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_661_inst_req_1;
      MUX_661_inst_ack_1<= update_ack(0);
      MUX_661_inst: SelectSplitProtocol generic map(name => "MUX_661_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_656_wire, y => type_cast_660_wire, sel => UGE_u2_u1_652_wire, z => col_to_be_replaced_2_662, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_673_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_673_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_673_inst:started:   inputs: " & " EQ_u2_u1_666_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_666_wire) & " type_cast_668_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_668_wire_constant) & " type_cast_672_wire = "& Convert_SLV_To_Hex_String(type_cast_672_wire));
          --
        end if; 
        if MUX_673_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUX_673_inst:finished:  outputs: " & " col_to_be_replaced_3_674= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_3_674));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_673_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_673_inst_req_0;
      MUX_673_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_673_inst_req_1;
      MUX_673_inst_ack_1<= update_ack(0);
      MUX_673_inst: SelectSplitProtocol generic map(name => "MUX_673_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_668_wire_constant, y => type_cast_672_wire, sel => EQ_u2_u1_666_wire, z => col_to_be_replaced_3_674, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator type_cast_646_inst flow-through 
    process(type_cast_646_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_646_inst:flowthrough inputs: " & " SUB_u2_u2_645_wire = "& Convert_SLV_To_Hex_String(SUB_u2_u2_645_wire) & " outputs:" & " type_cast_646_wire= "  & Convert_SLV_To_Hex_String(type_cast_646_wire));
      --
    end process; 
    -- interlock type_cast_646_inst
    process(SUB_u2_u2_645_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := SUB_u2_u2_645_wire(1 downto 0);
      type_cast_646_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_656_inst flow-through 
    process(type_cast_656_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_656_inst:flowthrough inputs: " & " SUB_u2_u2_655_wire = "& Convert_SLV_To_Hex_String(SUB_u2_u2_655_wire) & " outputs:" & " type_cast_656_wire= "  & Convert_SLV_To_Hex_String(type_cast_656_wire));
      --
    end process; 
    -- interlock type_cast_656_inst
    process(SUB_u2_u2_655_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := SUB_u2_u2_655_wire(1 downto 0);
      type_cast_656_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_660_inst flow-through 
    process(type_cast_660_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_660_inst:flowthrough inputs: " & " ADD_u2_u2_659_wire = "& Convert_SLV_To_Hex_String(ADD_u2_u2_659_wire) & " outputs:" & " type_cast_660_wire= "  & Convert_SLV_To_Hex_String(type_cast_660_wire));
      --
    end process; 
    -- interlock type_cast_660_inst
    process(ADD_u2_u2_659_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := ADD_u2_u2_659_wire(1 downto 0);
      type_cast_660_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_672_inst flow-through 
    process(type_cast_672_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_672_inst:flowthrough inputs: " & " ADD_u2_u2_671_wire = "& Convert_SLV_To_Hex_String(ADD_u2_u2_671_wire) & " outputs:" & " type_cast_672_wire= "  & Convert_SLV_To_Hex_String(type_cast_672_wire));
      --
    end process; 
    -- interlock type_cast_672_inst
    process(ADD_u2_u2_671_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := ADD_u2_u2_671_wire(1 downto 0);
      type_cast_672_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_683_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_683_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_683_inst:started:   inputs: " & " MUL_u16_u16_682_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_682_wire));
          --
        end if; 
        if type_cast_683_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_683_inst:finished:  outputs: " & " pp03_684= "  & Convert_SLV_To_Hex_String(pp03_684));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_683_inst_req_0;
      type_cast_683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_683_inst_req_1;
      type_cast_683_inst_ack_1<= rack(0);
      type_cast_683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_683_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_682_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp03_684,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_693_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_693_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_693_inst:started:   inputs: " & " MUL_u16_u16_692_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_692_wire));
          --
        end if; 
        if type_cast_693_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_693_inst:finished:  outputs: " & " pp13_694= "  & Convert_SLV_To_Hex_String(pp13_694));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_693_inst_req_0;
      type_cast_693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_693_inst_req_1;
      type_cast_693_inst_ack_1<= rack(0);
      type_cast_693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_692_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp13_694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_703_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_703_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_703_inst:started:   inputs: " & " MUL_u16_u16_702_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_702_wire));
          --
        end if; 
        if type_cast_703_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_703_inst:finished:  outputs: " & " pp23_704= "  & Convert_SLV_To_Hex_String(pp23_704));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_703_inst_req_0;
      type_cast_703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_703_inst_req_1;
      type_cast_703_inst_ack_1<= rack(0);
      type_cast_703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_702_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp23_704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_713_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_713_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_713_inst:started:   inputs: " & " MUL_u16_u16_712_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_712_wire));
          --
        end if; 
        if type_cast_713_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_713_inst:finished:  outputs: " & " pp33_714= "  & Convert_SLV_To_Hex_String(pp33_714));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_713_inst_req_0;
      type_cast_713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_713_inst_req_1;
      type_cast_713_inst_ack_1<= rack(0);
      type_cast_713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_712_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp33_714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_723_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_723_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_723_inst:started:   inputs: " & " MUL_u16_u16_722_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_722_wire));
          --
        end if; 
        if type_cast_723_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_723_inst:finished:  outputs: " & " pp02_724= "  & Convert_SLV_To_Hex_String(pp02_724));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_723_inst_req_0;
      type_cast_723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_723_inst_req_1;
      type_cast_723_inst_ack_1<= rack(0);
      type_cast_723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_722_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp02_724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_733_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_733_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_733_inst:started:   inputs: " & " MUL_u16_u16_732_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_732_wire));
          --
        end if; 
        if type_cast_733_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_733_inst:finished:  outputs: " & " pp12_734= "  & Convert_SLV_To_Hex_String(pp12_734));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_733_inst_req_0;
      type_cast_733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_733_inst_req_1;
      type_cast_733_inst_ack_1<= rack(0);
      type_cast_733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_732_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp12_734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_743_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_743_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_743_inst:started:   inputs: " & " MUL_u16_u16_742_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_742_wire));
          --
        end if; 
        if type_cast_743_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_743_inst:finished:  outputs: " & " pp22_744= "  & Convert_SLV_To_Hex_String(pp22_744));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_743_inst_req_0;
      type_cast_743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_743_inst_req_1;
      type_cast_743_inst_ack_1<= rack(0);
      type_cast_743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_742_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp22_744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_753_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_753_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_753_inst:started:   inputs: " & " MUL_u16_u16_752_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_752_wire));
          --
        end if; 
        if type_cast_753_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_753_inst:finished:  outputs: " & " pp32_754= "  & Convert_SLV_To_Hex_String(pp32_754));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_753_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_753_inst_req_0;
      type_cast_753_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_753_inst_req_1;
      type_cast_753_inst_ack_1<= rack(0);
      type_cast_753_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_753_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_752_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp32_754,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_763_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_763_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_763_inst:started:   inputs: " & " MUL_u16_u16_762_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_762_wire));
          --
        end if; 
        if type_cast_763_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_763_inst:finished:  outputs: " & " pp01_764= "  & Convert_SLV_To_Hex_String(pp01_764));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_762_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp01_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_773_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_773_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_773_inst:started:   inputs: " & " MUL_u16_u16_772_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_772_wire));
          --
        end if; 
        if type_cast_773_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_773_inst:finished:  outputs: " & " pp11_774= "  & Convert_SLV_To_Hex_String(pp11_774));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_773_inst_req_0;
      type_cast_773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_773_inst_req_1;
      type_cast_773_inst_ack_1<= rack(0);
      type_cast_773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_772_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp11_774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_783_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_783_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_783_inst:started:   inputs: " & " MUL_u16_u16_782_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_782_wire));
          --
        end if; 
        if type_cast_783_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_783_inst:finished:  outputs: " & " pp21_784= "  & Convert_SLV_To_Hex_String(pp21_784));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_783_inst_req_0;
      type_cast_783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_783_inst_req_1;
      type_cast_783_inst_ack_1<= rack(0);
      type_cast_783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_782_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp21_784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_793_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_793_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_793_inst:started:   inputs: " & " MUL_u16_u16_792_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_792_wire));
          --
        end if; 
        if type_cast_793_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_793_inst:finished:  outputs: " & " pp31_794= "  & Convert_SLV_To_Hex_String(pp31_794));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_792_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp31_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_803_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_803_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_803_inst:started:   inputs: " & " MUL_u16_u16_802_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_802_wire));
          --
        end if; 
        if type_cast_803_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_803_inst:finished:  outputs: " & " pp00_804= "  & Convert_SLV_To_Hex_String(pp00_804));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_803_inst_req_0;
      type_cast_803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_803_inst_req_1;
      type_cast_803_inst_ack_1<= rack(0);
      type_cast_803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_802_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp00_804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_813_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_813_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_813_inst:started:   inputs: " & " MUL_u16_u16_812_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_812_wire));
          --
        end if; 
        if type_cast_813_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_813_inst:finished:  outputs: " & " pp10_814= "  & Convert_SLV_To_Hex_String(pp10_814));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_813_inst_req_0;
      type_cast_813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_813_inst_req_1;
      type_cast_813_inst_ack_1<= rack(0);
      type_cast_813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_812_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp10_814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_823_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_823_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_823_inst:started:   inputs: " & " MUL_u16_u16_822_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_822_wire));
          --
        end if; 
        if type_cast_823_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_823_inst:finished:  outputs: " & " pp20_824= "  & Convert_SLV_To_Hex_String(pp20_824));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_823_inst_req_0;
      type_cast_823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_823_inst_req_1;
      type_cast_823_inst_ack_1<= rack(0);
      type_cast_823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_822_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp20_824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_833_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_833_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_833_inst:started:   inputs: " & " MUL_u16_u16_832_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_832_wire));
          --
        end if; 
        if type_cast_833_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_833_inst:finished:  outputs: " & " pp30_834= "  & Convert_SLV_To_Hex_String(pp30_834));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_833_inst_req_1;
      type_cast_833_inst_ack_1<= rack(0);
      type_cast_833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_832_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp30_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_839_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_839_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_839_inst:started:   inputs: " & " ADD_u16_u16_838_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_838_wire));
          --
        end if; 
        if type_cast_839_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_839_inst:finished:  outputs: " & " sum0_840= "  & Convert_SLV_To_Hex_String(sum0_840));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_839_inst_req_0;
      type_cast_839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_839_inst_req_1;
      type_cast_839_inst_ack_1<= rack(0);
      type_cast_839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_838_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum0_840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_845_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_845_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_845_inst:started:   inputs: " & " ADD_u16_u16_844_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_844_wire));
          --
        end if; 
        if type_cast_845_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_845_inst:finished:  outputs: " & " sum1_846= "  & Convert_SLV_To_Hex_String(sum1_846));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_845_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_845_inst_req_0;
      type_cast_845_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_845_inst_req_1;
      type_cast_845_inst_ack_1<= rack(0);
      type_cast_845_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_845_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_844_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum1_846,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_851_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_851_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_851_inst:started:   inputs: " & " ADD_u16_u16_850_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_850_wire));
          --
        end if; 
        if type_cast_851_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_851_inst:finished:  outputs: " & " sum2_852= "  & Convert_SLV_To_Hex_String(sum2_852));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_850_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum2_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_857_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_857_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_857_inst:started:   inputs: " & " ADD_u16_u16_856_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_856_wire));
          --
        end if; 
        if type_cast_857_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_857_inst:finished:  outputs: " & " sum3_858= "  & Convert_SLV_To_Hex_String(sum3_858));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_857_inst_req_0;
      type_cast_857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_857_inst_req_1;
      type_cast_857_inst_ack_1<= rack(0);
      type_cast_857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_856_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum3_858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_863_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_863_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_863_inst:started:   inputs: " & " ADD_u16_u16_862_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_862_wire));
          --
        end if; 
        if type_cast_863_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_863_inst:finished:  outputs: " & " sum4_864= "  & Convert_SLV_To_Hex_String(sum4_864));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_863_inst_req_1;
      type_cast_863_inst_ack_1<= rack(0);
      type_cast_863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_862_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum4_864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_869_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_869_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_869_inst:started:   inputs: " & " ADD_u16_u16_868_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_868_wire));
          --
        end if; 
        if type_cast_869_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_869_inst:finished:  outputs: " & " sum5_870= "  & Convert_SLV_To_Hex_String(sum5_870));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_869_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_869_inst_req_0;
      type_cast_869_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_869_inst_req_1;
      type_cast_869_inst_ack_1<= rack(0);
      type_cast_869_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_869_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_868_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum5_870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_875_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_875_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_875_inst:started:   inputs: " & " ADD_u16_u16_874_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_874_wire));
          --
        end if; 
        if type_cast_875_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_875_inst:finished:  outputs: " & " sum6_876= "  & Convert_SLV_To_Hex_String(sum6_876));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_875_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_875_inst_req_0;
      type_cast_875_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_875_inst_req_1;
      type_cast_875_inst_ack_1<= rack(0);
      type_cast_875_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_875_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_874_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum6_876,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_881_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_881_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_881_inst:started:   inputs: " & " ADD_u16_u16_880_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_880_wire));
          --
        end if; 
        if type_cast_881_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_881_inst:finished:  outputs: " & " sum7_882= "  & Convert_SLV_To_Hex_String(sum7_882));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_881_inst_req_0;
      type_cast_881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_881_inst_req_1;
      type_cast_881_inst_ack_1<= rack(0);
      type_cast_881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_880_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum7_882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_887_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_887_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_887_inst:started:   inputs: " & " ADD_u16_u16_886_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_886_wire));
          --
        end if; 
        if type_cast_887_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_887_inst:finished:  outputs: " & " sum10_888= "  & Convert_SLV_To_Hex_String(sum10_888));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_886_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum10_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_893_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_893_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_893_inst:started:   inputs: " & " ADD_u16_u16_892_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_892_wire));
          --
        end if; 
        if type_cast_893_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_893_inst:finished:  outputs: " & " sum11_894= "  & Convert_SLV_To_Hex_String(sum11_894));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_893_inst_req_0;
      type_cast_893_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_893_inst_req_1;
      type_cast_893_inst_ack_1<= rack(0);
      type_cast_893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_892_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum11_894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_899_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_899_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_899_inst:started:   inputs: " & " ADD_u16_u16_898_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_898_wire));
          --
        end if; 
        if type_cast_899_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_899_inst:finished:  outputs: " & " sum12_900= "  & Convert_SLV_To_Hex_String(sum12_900));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_899_inst_req_0;
      type_cast_899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_899_inst_req_1;
      type_cast_899_inst_ack_1<= rack(0);
      type_cast_899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_898_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum12_900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_905_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_905_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_905_inst:started:   inputs: " & " ADD_u16_u16_904_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_904_wire));
          --
        end if; 
        if type_cast_905_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_905_inst:finished:  outputs: " & " sum13_906= "  & Convert_SLV_To_Hex_String(sum13_906));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_904_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum13_906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_911_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_911_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_911_inst:started:   inputs: " & " ADD_u16_u16_910_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_910_wire));
          --
        end if; 
        if type_cast_911_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_911_inst:finished:  outputs: " & " sum20_912= "  & Convert_SLV_To_Hex_String(sum20_912));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_911_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_911_inst_req_0;
      type_cast_911_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_911_inst_req_1;
      type_cast_911_inst_ack_1<= rack(0);
      type_cast_911_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_911_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_910_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum20_912,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_917_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_917_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_917_inst:started:   inputs: " & " ADD_u16_u16_916_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_916_wire));
          --
        end if; 
        if type_cast_917_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_917_inst:finished:  outputs: " & " sum21_918= "  & Convert_SLV_To_Hex_String(sum21_918));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_917_inst_req_0;
      type_cast_917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_917_inst_req_1;
      type_cast_917_inst_ack_1<= rack(0);
      type_cast_917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_916_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum21_918,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_923_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_923_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_923_inst:started:   inputs: " & " ADD_u16_u16_922_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_922_wire));
          --
        end if; 
        if type_cast_923_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:type_cast_923_inst:finished:  outputs: " & " ofmap_pixel_buffer= "  & Convert_SLV_To_Hex_String(ofmap_pixel_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_922_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ofmap_pixel_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_678_addr_0 flow-through 
    process(array_obj_ref_678_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_addr_0:flowthrough  inputs: " & " array_obj_ref_678_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_678_root_address) & "outputs: " & " array_obj_ref_678_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_678_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_678_addr_0
    process(array_obj_ref_678_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_678_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_678_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_678_gather_scatter flow-through 
    process(array_obj_ref_678_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_gather_scatter:flowthrough  inputs: " & " array_obj_ref_678_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_678_data_0) & "outputs: " & " array_obj_ref_678_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_678_wire));
      --
    end process; 
    -- equivalence array_obj_ref_678_gather_scatter
    process(array_obj_ref_678_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_678_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_678_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_678_index_1_rename flow-through 
    process(R_col_to_be_replaced_677_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_677_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_677_resized) & "outputs: " & " R_col_to_be_replaced_677_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_677_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_678_index_1_rename
    process(R_col_to_be_replaced_677_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_677_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_677_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_678_index_1_resize flow-through 
    process(R_col_to_be_replaced_677_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_677_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_677_resized));
      --
    end process; 
    -- equivalence array_obj_ref_678_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_677_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_678_root_address_inst flow-through 
    process(array_obj_ref_678_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_root_address_inst:flowthrough  inputs: " & " array_obj_ref_678_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_678_final_offset) & "outputs: " & " array_obj_ref_678_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_678_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_678_root_address_inst
    process(array_obj_ref_678_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_678_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_678_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_681_gather_scatter flow-through 
    process(array_obj_ref_681_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_681_gather_scatter:flowthrough  inputs: " & " array_obj_ref_681_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_681_data_0) & "outputs: " & " array_obj_ref_681_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_681_wire));
      --
    end process; 
    -- equivalence array_obj_ref_681_gather_scatter
    process(array_obj_ref_681_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_681_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_681_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_688_addr_0 flow-through 
    process(array_obj_ref_688_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_addr_0:flowthrough  inputs: " & " array_obj_ref_688_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_688_root_address) & "outputs: " & " array_obj_ref_688_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_688_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_688_addr_0
    process(array_obj_ref_688_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_688_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_688_gather_scatter flow-through 
    process(array_obj_ref_688_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_gather_scatter:flowthrough  inputs: " & " array_obj_ref_688_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_688_data_0) & "outputs: " & " array_obj_ref_688_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_688_wire));
      --
    end process; 
    -- equivalence array_obj_ref_688_gather_scatter
    process(array_obj_ref_688_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_688_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_688_index_1_rename flow-through 
    process(R_col_to_be_replaced_687_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_687_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_687_resized) & "outputs: " & " R_col_to_be_replaced_687_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_687_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_688_index_1_rename
    process(R_col_to_be_replaced_687_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_687_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_687_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_688_index_1_resize flow-through 
    process(R_col_to_be_replaced_687_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_687_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_687_resized));
      --
    end process; 
    -- equivalence array_obj_ref_688_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_687_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_688_root_address_inst flow-through 
    process(array_obj_ref_688_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_root_address_inst:flowthrough  inputs: " & " array_obj_ref_688_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_688_final_offset) & "outputs: " & " array_obj_ref_688_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_688_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_688_root_address_inst
    process(array_obj_ref_688_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_688_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_691_gather_scatter flow-through 
    process(array_obj_ref_691_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_691_gather_scatter:flowthrough  inputs: " & " array_obj_ref_691_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_691_data_0) & "outputs: " & " array_obj_ref_691_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_691_wire));
      --
    end process; 
    -- equivalence array_obj_ref_691_gather_scatter
    process(array_obj_ref_691_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_691_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_691_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_698_addr_0 flow-through 
    process(array_obj_ref_698_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_addr_0:flowthrough  inputs: " & " array_obj_ref_698_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_698_root_address) & "outputs: " & " array_obj_ref_698_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_698_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_698_addr_0
    process(array_obj_ref_698_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_698_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_698_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_698_gather_scatter flow-through 
    process(array_obj_ref_698_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_gather_scatter:flowthrough  inputs: " & " array_obj_ref_698_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_698_data_0) & "outputs: " & " array_obj_ref_698_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_698_wire));
      --
    end process; 
    -- equivalence array_obj_ref_698_gather_scatter
    process(array_obj_ref_698_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_698_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_698_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_698_index_1_rename flow-through 
    process(R_col_to_be_replaced_697_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_697_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_697_resized) & "outputs: " & " R_col_to_be_replaced_697_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_697_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_698_index_1_rename
    process(R_col_to_be_replaced_697_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_697_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_697_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_698_index_1_resize flow-through 
    process(R_col_to_be_replaced_697_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_697_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_697_resized));
      --
    end process; 
    -- equivalence array_obj_ref_698_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_697_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_698_root_address_inst flow-through 
    process(array_obj_ref_698_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_root_address_inst:flowthrough  inputs: " & " array_obj_ref_698_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_698_final_offset) & "outputs: " & " array_obj_ref_698_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_698_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_698_root_address_inst
    process(array_obj_ref_698_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_698_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_698_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_701_gather_scatter flow-through 
    process(array_obj_ref_701_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_701_gather_scatter:flowthrough  inputs: " & " array_obj_ref_701_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_701_data_0) & "outputs: " & " array_obj_ref_701_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_701_wire));
      --
    end process; 
    -- equivalence array_obj_ref_701_gather_scatter
    process(array_obj_ref_701_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_701_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_701_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_708_addr_0 flow-through 
    process(array_obj_ref_708_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_addr_0:flowthrough  inputs: " & " array_obj_ref_708_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_708_root_address) & "outputs: " & " array_obj_ref_708_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_708_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_708_addr_0
    process(array_obj_ref_708_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_708_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_708_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_708_gather_scatter flow-through 
    process(array_obj_ref_708_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_gather_scatter:flowthrough  inputs: " & " array_obj_ref_708_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_708_data_0) & "outputs: " & " array_obj_ref_708_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_708_wire));
      --
    end process; 
    -- equivalence array_obj_ref_708_gather_scatter
    process(array_obj_ref_708_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_708_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_708_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_708_index_1_rename flow-through 
    process(R_col_to_be_replaced_707_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_707_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_707_resized) & "outputs: " & " R_col_to_be_replaced_707_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_707_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_708_index_1_rename
    process(R_col_to_be_replaced_707_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_707_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_707_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_708_index_1_resize flow-through 
    process(R_col_to_be_replaced_707_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_707_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_707_resized));
      --
    end process; 
    -- equivalence array_obj_ref_708_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_707_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_708_root_address_inst flow-through 
    process(array_obj_ref_708_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_root_address_inst:flowthrough  inputs: " & " array_obj_ref_708_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_708_final_offset) & "outputs: " & " array_obj_ref_708_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_708_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_708_root_address_inst
    process(array_obj_ref_708_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_708_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_708_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_711_gather_scatter flow-through 
    process(array_obj_ref_711_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_711_gather_scatter:flowthrough  inputs: " & " array_obj_ref_711_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_711_data_0) & "outputs: " & " array_obj_ref_711_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_711_wire));
      --
    end process; 
    -- equivalence array_obj_ref_711_gather_scatter
    process(array_obj_ref_711_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_711_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_711_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_718_addr_0 flow-through 
    process(array_obj_ref_718_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_addr_0:flowthrough  inputs: " & " array_obj_ref_718_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_718_root_address) & "outputs: " & " array_obj_ref_718_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_718_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_718_addr_0
    process(array_obj_ref_718_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_718_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_718_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_718_gather_scatter flow-through 
    process(array_obj_ref_718_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_gather_scatter:flowthrough  inputs: " & " array_obj_ref_718_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_718_data_0) & "outputs: " & " array_obj_ref_718_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_718_wire));
      --
    end process; 
    -- equivalence array_obj_ref_718_gather_scatter
    process(array_obj_ref_718_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_718_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_718_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_718_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_717_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_717_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_717_resized) & "outputs: " & " R_col_to_be_replaced_1_717_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_717_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_718_index_1_rename
    process(R_col_to_be_replaced_1_717_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_717_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_717_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_718_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_717_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_648 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_648) & "outputs: " & " R_col_to_be_replaced_1_717_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_717_resized));
      --
    end process; 
    -- equivalence array_obj_ref_718_index_1_resize
    process(col_to_be_replaced_1_648) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_648;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_717_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_718_root_address_inst flow-through 
    process(array_obj_ref_718_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_root_address_inst:flowthrough  inputs: " & " array_obj_ref_718_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_718_final_offset) & "outputs: " & " array_obj_ref_718_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_718_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_718_root_address_inst
    process(array_obj_ref_718_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_718_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_718_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_721_gather_scatter flow-through 
    process(array_obj_ref_721_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_721_gather_scatter:flowthrough  inputs: " & " array_obj_ref_721_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_721_data_0) & "outputs: " & " array_obj_ref_721_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_721_wire));
      --
    end process; 
    -- equivalence array_obj_ref_721_gather_scatter
    process(array_obj_ref_721_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_721_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_721_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_728_addr_0 flow-through 
    process(array_obj_ref_728_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_addr_0:flowthrough  inputs: " & " array_obj_ref_728_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_728_root_address) & "outputs: " & " array_obj_ref_728_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_728_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_728_addr_0
    process(array_obj_ref_728_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_728_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_728_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_728_gather_scatter flow-through 
    process(array_obj_ref_728_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_gather_scatter:flowthrough  inputs: " & " array_obj_ref_728_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_728_data_0) & "outputs: " & " array_obj_ref_728_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_728_wire));
      --
    end process; 
    -- equivalence array_obj_ref_728_gather_scatter
    process(array_obj_ref_728_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_728_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_728_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_728_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_727_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_727_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_727_resized) & "outputs: " & " R_col_to_be_replaced_1_727_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_727_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_728_index_1_rename
    process(R_col_to_be_replaced_1_727_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_727_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_727_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_728_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_727_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_648 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_648) & "outputs: " & " R_col_to_be_replaced_1_727_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_727_resized));
      --
    end process; 
    -- equivalence array_obj_ref_728_index_1_resize
    process(col_to_be_replaced_1_648) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_648;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_727_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_728_root_address_inst flow-through 
    process(array_obj_ref_728_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_root_address_inst:flowthrough  inputs: " & " array_obj_ref_728_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_728_final_offset) & "outputs: " & " array_obj_ref_728_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_728_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_728_root_address_inst
    process(array_obj_ref_728_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_728_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_728_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_731_gather_scatter flow-through 
    process(array_obj_ref_731_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_731_gather_scatter:flowthrough  inputs: " & " array_obj_ref_731_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_731_data_0) & "outputs: " & " array_obj_ref_731_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_731_wire));
      --
    end process; 
    -- equivalence array_obj_ref_731_gather_scatter
    process(array_obj_ref_731_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_731_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_731_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_738_addr_0 flow-through 
    process(array_obj_ref_738_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_addr_0:flowthrough  inputs: " & " array_obj_ref_738_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_738_root_address) & "outputs: " & " array_obj_ref_738_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_738_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_738_addr_0
    process(array_obj_ref_738_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_738_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_738_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_738_gather_scatter flow-through 
    process(array_obj_ref_738_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_gather_scatter:flowthrough  inputs: " & " array_obj_ref_738_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_738_data_0) & "outputs: " & " array_obj_ref_738_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_738_wire));
      --
    end process; 
    -- equivalence array_obj_ref_738_gather_scatter
    process(array_obj_ref_738_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_738_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_738_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_738_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_737_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_737_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_737_resized) & "outputs: " & " R_col_to_be_replaced_1_737_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_737_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_738_index_1_rename
    process(R_col_to_be_replaced_1_737_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_737_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_737_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_738_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_737_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_648 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_648) & "outputs: " & " R_col_to_be_replaced_1_737_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_737_resized));
      --
    end process; 
    -- equivalence array_obj_ref_738_index_1_resize
    process(col_to_be_replaced_1_648) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_648;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_737_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_738_root_address_inst flow-through 
    process(array_obj_ref_738_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_root_address_inst:flowthrough  inputs: " & " array_obj_ref_738_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_738_final_offset) & "outputs: " & " array_obj_ref_738_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_738_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_738_root_address_inst
    process(array_obj_ref_738_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_738_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_738_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_741_gather_scatter flow-through 
    process(array_obj_ref_741_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_741_gather_scatter:flowthrough  inputs: " & " array_obj_ref_741_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_741_data_0) & "outputs: " & " array_obj_ref_741_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_741_wire));
      --
    end process; 
    -- equivalence array_obj_ref_741_gather_scatter
    process(array_obj_ref_741_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_741_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_741_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_748_addr_0 flow-through 
    process(array_obj_ref_748_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_addr_0:flowthrough  inputs: " & " array_obj_ref_748_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_748_root_address) & "outputs: " & " array_obj_ref_748_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_748_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_748_addr_0
    process(array_obj_ref_748_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_748_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_748_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_748_gather_scatter flow-through 
    process(array_obj_ref_748_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_gather_scatter:flowthrough  inputs: " & " array_obj_ref_748_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_748_data_0) & "outputs: " & " array_obj_ref_748_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_748_wire));
      --
    end process; 
    -- equivalence array_obj_ref_748_gather_scatter
    process(array_obj_ref_748_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_748_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_748_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_748_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_747_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_747_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_747_resized) & "outputs: " & " R_col_to_be_replaced_1_747_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_747_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_748_index_1_rename
    process(R_col_to_be_replaced_1_747_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_747_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_747_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_748_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_747_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_648 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_648) & "outputs: " & " R_col_to_be_replaced_1_747_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_747_resized));
      --
    end process; 
    -- equivalence array_obj_ref_748_index_1_resize
    process(col_to_be_replaced_1_648) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_648;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_747_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_748_root_address_inst flow-through 
    process(array_obj_ref_748_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_root_address_inst:flowthrough  inputs: " & " array_obj_ref_748_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_748_final_offset) & "outputs: " & " array_obj_ref_748_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_748_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_748_root_address_inst
    process(array_obj_ref_748_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_748_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_748_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_751_gather_scatter flow-through 
    process(array_obj_ref_751_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_751_gather_scatter:flowthrough  inputs: " & " array_obj_ref_751_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_751_data_0) & "outputs: " & " array_obj_ref_751_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_751_wire));
      --
    end process; 
    -- equivalence array_obj_ref_751_gather_scatter
    process(array_obj_ref_751_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_751_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_751_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_758_addr_0 flow-through 
    process(array_obj_ref_758_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_addr_0:flowthrough  inputs: " & " array_obj_ref_758_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_758_root_address) & "outputs: " & " array_obj_ref_758_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_758_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_758_addr_0
    process(array_obj_ref_758_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_758_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_758_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_758_gather_scatter flow-through 
    process(array_obj_ref_758_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_gather_scatter:flowthrough  inputs: " & " array_obj_ref_758_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_758_data_0) & "outputs: " & " array_obj_ref_758_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_758_wire));
      --
    end process; 
    -- equivalence array_obj_ref_758_gather_scatter
    process(array_obj_ref_758_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_758_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_758_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_758_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_757_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_757_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_757_resized) & "outputs: " & " R_col_to_be_replaced_2_757_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_757_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_758_index_1_rename
    process(R_col_to_be_replaced_2_757_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_757_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_757_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_758_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_757_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_662 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_662) & "outputs: " & " R_col_to_be_replaced_2_757_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_757_resized));
      --
    end process; 
    -- equivalence array_obj_ref_758_index_1_resize
    process(col_to_be_replaced_2_662) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_662;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_757_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_758_root_address_inst flow-through 
    process(array_obj_ref_758_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_root_address_inst:flowthrough  inputs: " & " array_obj_ref_758_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_758_final_offset) & "outputs: " & " array_obj_ref_758_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_758_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_758_root_address_inst
    process(array_obj_ref_758_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_758_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_758_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_761_gather_scatter flow-through 
    process(array_obj_ref_761_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_761_gather_scatter:flowthrough  inputs: " & " array_obj_ref_761_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_761_data_0) & "outputs: " & " array_obj_ref_761_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_761_wire));
      --
    end process; 
    -- equivalence array_obj_ref_761_gather_scatter
    process(array_obj_ref_761_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_761_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_761_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_768_addr_0 flow-through 
    process(array_obj_ref_768_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_addr_0:flowthrough  inputs: " & " array_obj_ref_768_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_768_root_address) & "outputs: " & " array_obj_ref_768_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_768_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_768_addr_0
    process(array_obj_ref_768_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_768_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_768_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_768_gather_scatter flow-through 
    process(array_obj_ref_768_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_gather_scatter:flowthrough  inputs: " & " array_obj_ref_768_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_768_data_0) & "outputs: " & " array_obj_ref_768_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_768_wire));
      --
    end process; 
    -- equivalence array_obj_ref_768_gather_scatter
    process(array_obj_ref_768_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_768_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_768_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_768_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_767_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_767_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_767_resized) & "outputs: " & " R_col_to_be_replaced_2_767_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_767_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_768_index_1_rename
    process(R_col_to_be_replaced_2_767_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_767_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_767_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_768_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_767_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_662 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_662) & "outputs: " & " R_col_to_be_replaced_2_767_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_767_resized));
      --
    end process; 
    -- equivalence array_obj_ref_768_index_1_resize
    process(col_to_be_replaced_2_662) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_662;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_767_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_768_root_address_inst flow-through 
    process(array_obj_ref_768_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_root_address_inst:flowthrough  inputs: " & " array_obj_ref_768_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_768_final_offset) & "outputs: " & " array_obj_ref_768_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_768_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_768_root_address_inst
    process(array_obj_ref_768_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_768_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_768_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_771_gather_scatter flow-through 
    process(array_obj_ref_771_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_771_gather_scatter:flowthrough  inputs: " & " array_obj_ref_771_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_771_data_0) & "outputs: " & " array_obj_ref_771_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_771_wire));
      --
    end process; 
    -- equivalence array_obj_ref_771_gather_scatter
    process(array_obj_ref_771_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_771_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_771_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_778_addr_0 flow-through 
    process(array_obj_ref_778_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_addr_0:flowthrough  inputs: " & " array_obj_ref_778_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_778_root_address) & "outputs: " & " array_obj_ref_778_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_778_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_778_addr_0
    process(array_obj_ref_778_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_778_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_778_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_778_gather_scatter flow-through 
    process(array_obj_ref_778_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_gather_scatter:flowthrough  inputs: " & " array_obj_ref_778_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_778_data_0) & "outputs: " & " array_obj_ref_778_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_778_wire));
      --
    end process; 
    -- equivalence array_obj_ref_778_gather_scatter
    process(array_obj_ref_778_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_778_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_778_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_778_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_777_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_777_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_777_resized) & "outputs: " & " R_col_to_be_replaced_2_777_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_777_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_778_index_1_rename
    process(R_col_to_be_replaced_2_777_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_777_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_777_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_778_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_777_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_662 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_662) & "outputs: " & " R_col_to_be_replaced_2_777_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_777_resized));
      --
    end process; 
    -- equivalence array_obj_ref_778_index_1_resize
    process(col_to_be_replaced_2_662) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_662;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_777_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_778_root_address_inst flow-through 
    process(array_obj_ref_778_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_root_address_inst:flowthrough  inputs: " & " array_obj_ref_778_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_778_final_offset) & "outputs: " & " array_obj_ref_778_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_778_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_778_root_address_inst
    process(array_obj_ref_778_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_778_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_778_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_781_gather_scatter flow-through 
    process(array_obj_ref_781_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_781_gather_scatter:flowthrough  inputs: " & " array_obj_ref_781_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_781_data_0) & "outputs: " & " array_obj_ref_781_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_781_wire));
      --
    end process; 
    -- equivalence array_obj_ref_781_gather_scatter
    process(array_obj_ref_781_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_781_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_781_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_788_addr_0 flow-through 
    process(array_obj_ref_788_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_addr_0:flowthrough  inputs: " & " array_obj_ref_788_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_788_root_address) & "outputs: " & " array_obj_ref_788_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_788_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_788_addr_0
    process(array_obj_ref_788_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_788_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_788_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_788_gather_scatter flow-through 
    process(array_obj_ref_788_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_gather_scatter:flowthrough  inputs: " & " array_obj_ref_788_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_788_data_0) & "outputs: " & " array_obj_ref_788_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_788_wire));
      --
    end process; 
    -- equivalence array_obj_ref_788_gather_scatter
    process(array_obj_ref_788_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_788_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_788_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_788_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_787_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_787_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_787_resized) & "outputs: " & " R_col_to_be_replaced_2_787_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_787_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_788_index_1_rename
    process(R_col_to_be_replaced_2_787_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_787_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_787_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_788_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_787_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_662 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_662) & "outputs: " & " R_col_to_be_replaced_2_787_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_787_resized));
      --
    end process; 
    -- equivalence array_obj_ref_788_index_1_resize
    process(col_to_be_replaced_2_662) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_662;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_787_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_788_root_address_inst flow-through 
    process(array_obj_ref_788_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_root_address_inst:flowthrough  inputs: " & " array_obj_ref_788_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_788_final_offset) & "outputs: " & " array_obj_ref_788_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_788_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_788_root_address_inst
    process(array_obj_ref_788_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_788_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_788_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_791_gather_scatter flow-through 
    process(array_obj_ref_791_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_791_gather_scatter:flowthrough  inputs: " & " array_obj_ref_791_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_791_data_0) & "outputs: " & " array_obj_ref_791_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_791_wire));
      --
    end process; 
    -- equivalence array_obj_ref_791_gather_scatter
    process(array_obj_ref_791_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_791_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_791_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_798_addr_0 flow-through 
    process(array_obj_ref_798_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_addr_0:flowthrough  inputs: " & " array_obj_ref_798_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_798_root_address) & "outputs: " & " array_obj_ref_798_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_798_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_798_addr_0
    process(array_obj_ref_798_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_798_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_798_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_798_gather_scatter flow-through 
    process(array_obj_ref_798_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_gather_scatter:flowthrough  inputs: " & " array_obj_ref_798_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_798_data_0) & "outputs: " & " array_obj_ref_798_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_798_wire));
      --
    end process; 
    -- equivalence array_obj_ref_798_gather_scatter
    process(array_obj_ref_798_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_798_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_798_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_798_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_797_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_797_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_797_resized) & "outputs: " & " R_col_to_be_replaced_3_797_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_797_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_798_index_1_rename
    process(R_col_to_be_replaced_3_797_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_797_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_797_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_798_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_797_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_674 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_674) & "outputs: " & " R_col_to_be_replaced_3_797_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_797_resized));
      --
    end process; 
    -- equivalence array_obj_ref_798_index_1_resize
    process(col_to_be_replaced_3_674) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_674;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_797_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_798_root_address_inst flow-through 
    process(array_obj_ref_798_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_root_address_inst:flowthrough  inputs: " & " array_obj_ref_798_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_798_final_offset) & "outputs: " & " array_obj_ref_798_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_798_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_798_root_address_inst
    process(array_obj_ref_798_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_798_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_798_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_801_gather_scatter flow-through 
    process(array_obj_ref_801_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_801_gather_scatter:flowthrough  inputs: " & " array_obj_ref_801_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_801_data_0) & "outputs: " & " array_obj_ref_801_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_801_wire));
      --
    end process; 
    -- equivalence array_obj_ref_801_gather_scatter
    process(array_obj_ref_801_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_801_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_801_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_808_addr_0 flow-through 
    process(array_obj_ref_808_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_addr_0:flowthrough  inputs: " & " array_obj_ref_808_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_808_root_address) & "outputs: " & " array_obj_ref_808_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_808_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_808_addr_0
    process(array_obj_ref_808_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_808_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_808_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_808_gather_scatter flow-through 
    process(array_obj_ref_808_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_gather_scatter:flowthrough  inputs: " & " array_obj_ref_808_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_808_data_0) & "outputs: " & " array_obj_ref_808_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_808_wire));
      --
    end process; 
    -- equivalence array_obj_ref_808_gather_scatter
    process(array_obj_ref_808_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_808_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_808_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_808_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_807_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_807_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_807_resized) & "outputs: " & " R_col_to_be_replaced_3_807_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_807_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_808_index_1_rename
    process(R_col_to_be_replaced_3_807_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_807_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_807_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_808_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_807_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_674 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_674) & "outputs: " & " R_col_to_be_replaced_3_807_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_807_resized));
      --
    end process; 
    -- equivalence array_obj_ref_808_index_1_resize
    process(col_to_be_replaced_3_674) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_674;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_807_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_808_root_address_inst flow-through 
    process(array_obj_ref_808_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_root_address_inst:flowthrough  inputs: " & " array_obj_ref_808_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_808_final_offset) & "outputs: " & " array_obj_ref_808_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_808_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_808_root_address_inst
    process(array_obj_ref_808_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_808_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_808_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_811_gather_scatter flow-through 
    process(array_obj_ref_811_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_811_gather_scatter:flowthrough  inputs: " & " array_obj_ref_811_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_811_data_0) & "outputs: " & " array_obj_ref_811_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_811_wire));
      --
    end process; 
    -- equivalence array_obj_ref_811_gather_scatter
    process(array_obj_ref_811_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_811_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_811_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_818_addr_0 flow-through 
    process(array_obj_ref_818_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_addr_0:flowthrough  inputs: " & " array_obj_ref_818_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_818_root_address) & "outputs: " & " array_obj_ref_818_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_818_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_818_addr_0
    process(array_obj_ref_818_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_818_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_818_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_818_gather_scatter flow-through 
    process(array_obj_ref_818_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_gather_scatter:flowthrough  inputs: " & " array_obj_ref_818_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_818_data_0) & "outputs: " & " array_obj_ref_818_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_818_wire));
      --
    end process; 
    -- equivalence array_obj_ref_818_gather_scatter
    process(array_obj_ref_818_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_818_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_818_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_818_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_817_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_817_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_817_resized) & "outputs: " & " R_col_to_be_replaced_3_817_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_817_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_818_index_1_rename
    process(R_col_to_be_replaced_3_817_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_817_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_817_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_818_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_817_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_674 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_674) & "outputs: " & " R_col_to_be_replaced_3_817_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_817_resized));
      --
    end process; 
    -- equivalence array_obj_ref_818_index_1_resize
    process(col_to_be_replaced_3_674) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_674;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_817_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_818_root_address_inst flow-through 
    process(array_obj_ref_818_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_root_address_inst:flowthrough  inputs: " & " array_obj_ref_818_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_818_final_offset) & "outputs: " & " array_obj_ref_818_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_818_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_818_root_address_inst
    process(array_obj_ref_818_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_818_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_818_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_821_gather_scatter flow-through 
    process(array_obj_ref_821_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_821_gather_scatter:flowthrough  inputs: " & " array_obj_ref_821_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_821_data_0) & "outputs: " & " array_obj_ref_821_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_821_wire));
      --
    end process; 
    -- equivalence array_obj_ref_821_gather_scatter
    process(array_obj_ref_821_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_821_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_821_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_828_addr_0 flow-through 
    process(array_obj_ref_828_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_addr_0:flowthrough  inputs: " & " array_obj_ref_828_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_828_root_address) & "outputs: " & " array_obj_ref_828_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_828_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_828_addr_0
    process(array_obj_ref_828_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_828_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_828_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_828_gather_scatter flow-through 
    process(array_obj_ref_828_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_gather_scatter:flowthrough  inputs: " & " array_obj_ref_828_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_828_data_0) & "outputs: " & " array_obj_ref_828_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_828_wire));
      --
    end process; 
    -- equivalence array_obj_ref_828_gather_scatter
    process(array_obj_ref_828_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_828_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_828_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_828_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_827_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_827_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_827_resized) & "outputs: " & " R_col_to_be_replaced_3_827_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_827_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_828_index_1_rename
    process(R_col_to_be_replaced_3_827_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_827_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_827_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_828_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_827_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_674 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_674) & "outputs: " & " R_col_to_be_replaced_3_827_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_827_resized));
      --
    end process; 
    -- equivalence array_obj_ref_828_index_1_resize
    process(col_to_be_replaced_3_674) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_674;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_827_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_828_root_address_inst flow-through 
    process(array_obj_ref_828_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_root_address_inst:flowthrough  inputs: " & " array_obj_ref_828_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_828_final_offset) & "outputs: " & " array_obj_ref_828_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_828_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_828_root_address_inst
    process(array_obj_ref_828_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_828_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_828_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_831_gather_scatter flow-through 
    process(array_obj_ref_831_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_831_gather_scatter:flowthrough  inputs: " & " array_obj_ref_831_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_831_data_0) & "outputs: " & " array_obj_ref_831_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_831_wire));
      --
    end process; 
    -- equivalence array_obj_ref_831_gather_scatter
    process(array_obj_ref_831_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_831_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_831_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u16_u16_838_inst flow-through 
    process(ADD_u16_u16_838_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_838_inst:flowthrough inputs: " & " pp00_804 = "& Convert_SLV_To_Hex_String(pp00_804) & " pp01_764 = "& Convert_SLV_To_Hex_String(pp01_764) & " outputs:" & " ADD_u16_u16_838_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_838_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_838_inst
    process(pp00_804, pp01_764) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp00_804, pp01_764, tmp_var);
      ADD_u16_u16_838_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_844_inst flow-through 
    process(ADD_u16_u16_844_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_844_inst:flowthrough inputs: " & " pp02_724 = "& Convert_SLV_To_Hex_String(pp02_724) & " pp03_684 = "& Convert_SLV_To_Hex_String(pp03_684) & " outputs:" & " ADD_u16_u16_844_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_844_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_844_inst
    process(pp02_724, pp03_684) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp02_724, pp03_684, tmp_var);
      ADD_u16_u16_844_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_850_inst flow-through 
    process(ADD_u16_u16_850_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_850_inst:flowthrough inputs: " & " pp10_814 = "& Convert_SLV_To_Hex_String(pp10_814) & " pp11_774 = "& Convert_SLV_To_Hex_String(pp11_774) & " outputs:" & " ADD_u16_u16_850_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_850_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_850_inst
    process(pp10_814, pp11_774) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp10_814, pp11_774, tmp_var);
      ADD_u16_u16_850_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_856_inst flow-through 
    process(ADD_u16_u16_856_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_856_inst:flowthrough inputs: " & " pp12_734 = "& Convert_SLV_To_Hex_String(pp12_734) & " pp13_694 = "& Convert_SLV_To_Hex_String(pp13_694) & " outputs:" & " ADD_u16_u16_856_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_856_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_856_inst
    process(pp12_734, pp13_694) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp12_734, pp13_694, tmp_var);
      ADD_u16_u16_856_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_862_inst flow-through 
    process(ADD_u16_u16_862_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_862_inst:flowthrough inputs: " & " pp20_824 = "& Convert_SLV_To_Hex_String(pp20_824) & " pp21_784 = "& Convert_SLV_To_Hex_String(pp21_784) & " outputs:" & " ADD_u16_u16_862_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_862_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_862_inst
    process(pp20_824, pp21_784) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp20_824, pp21_784, tmp_var);
      ADD_u16_u16_862_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_868_inst flow-through 
    process(ADD_u16_u16_868_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_868_inst:flowthrough inputs: " & " pp22_744 = "& Convert_SLV_To_Hex_String(pp22_744) & " pp23_704 = "& Convert_SLV_To_Hex_String(pp23_704) & " outputs:" & " ADD_u16_u16_868_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_868_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_868_inst
    process(pp22_744, pp23_704) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp22_744, pp23_704, tmp_var);
      ADD_u16_u16_868_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_874_inst flow-through 
    process(ADD_u16_u16_874_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_874_inst:flowthrough inputs: " & " pp30_834 = "& Convert_SLV_To_Hex_String(pp30_834) & " pp31_794 = "& Convert_SLV_To_Hex_String(pp31_794) & " outputs:" & " ADD_u16_u16_874_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_874_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_874_inst
    process(pp30_834, pp31_794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp30_834, pp31_794, tmp_var);
      ADD_u16_u16_874_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_880_inst flow-through 
    process(ADD_u16_u16_880_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_880_inst:flowthrough inputs: " & " pp32_754 = "& Convert_SLV_To_Hex_String(pp32_754) & " pp33_714 = "& Convert_SLV_To_Hex_String(pp33_714) & " outputs:" & " ADD_u16_u16_880_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_880_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_880_inst
    process(pp32_754, pp33_714) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp32_754, pp33_714, tmp_var);
      ADD_u16_u16_880_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_886_inst flow-through 
    process(ADD_u16_u16_886_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_886_inst:flowthrough inputs: " & " sum0_840 = "& Convert_SLV_To_Hex_String(sum0_840) & " sum1_846 = "& Convert_SLV_To_Hex_String(sum1_846) & " outputs:" & " ADD_u16_u16_886_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_886_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_886_inst
    process(sum0_840, sum1_846) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum0_840, sum1_846, tmp_var);
      ADD_u16_u16_886_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_892_inst flow-through 
    process(ADD_u16_u16_892_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_892_inst:flowthrough inputs: " & " sum2_852 = "& Convert_SLV_To_Hex_String(sum2_852) & " sum3_858 = "& Convert_SLV_To_Hex_String(sum3_858) & " outputs:" & " ADD_u16_u16_892_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_892_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_892_inst
    process(sum2_852, sum3_858) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum2_852, sum3_858, tmp_var);
      ADD_u16_u16_892_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_898_inst flow-through 
    process(ADD_u16_u16_898_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_898_inst:flowthrough inputs: " & " sum4_864 = "& Convert_SLV_To_Hex_String(sum4_864) & " sum5_870 = "& Convert_SLV_To_Hex_String(sum5_870) & " outputs:" & " ADD_u16_u16_898_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_898_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_898_inst
    process(sum4_864, sum5_870) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum4_864, sum5_870, tmp_var);
      ADD_u16_u16_898_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_904_inst flow-through 
    process(ADD_u16_u16_904_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_904_inst:flowthrough inputs: " & " sum6_876 = "& Convert_SLV_To_Hex_String(sum6_876) & " sum7_882 = "& Convert_SLV_To_Hex_String(sum7_882) & " outputs:" & " ADD_u16_u16_904_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_904_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_904_inst
    process(sum6_876, sum7_882) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum6_876, sum7_882, tmp_var);
      ADD_u16_u16_904_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_910_inst flow-through 
    process(ADD_u16_u16_910_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_910_inst:flowthrough inputs: " & " sum10_888 = "& Convert_SLV_To_Hex_String(sum10_888) & " sum11_894 = "& Convert_SLV_To_Hex_String(sum11_894) & " outputs:" & " ADD_u16_u16_910_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_910_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_910_inst
    process(sum10_888, sum11_894) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum10_888, sum11_894, tmp_var);
      ADD_u16_u16_910_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_916_inst flow-through 
    process(ADD_u16_u16_916_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_916_inst:flowthrough inputs: " & " sum12_900 = "& Convert_SLV_To_Hex_String(sum12_900) & " sum13_906 = "& Convert_SLV_To_Hex_String(sum13_906) & " outputs:" & " ADD_u16_u16_916_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_916_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_916_inst
    process(sum12_900, sum13_906) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum12_900, sum13_906, tmp_var);
      ADD_u16_u16_916_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_922_inst flow-through 
    process(ADD_u16_u16_922_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u16_u16_922_inst:flowthrough inputs: " & " sum20_912 = "& Convert_SLV_To_Hex_String(sum20_912) & " sum21_918 = "& Convert_SLV_To_Hex_String(sum21_918) & " outputs:" & " ADD_u16_u16_922_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_922_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_922_inst
    process(sum20_912, sum21_918) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum20_912, sum21_918, tmp_var);
      ADD_u16_u16_922_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u2_u2_659_inst flow-through 
    process(ADD_u2_u2_659_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u2_u2_659_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_658_wire_constant = "& Convert_SLV_To_Hex_String(konst_658_wire_constant) & " outputs:" & " ADD_u2_u2_659_wire= "  & Convert_SLV_To_Hex_String(ADD_u2_u2_659_wire));
      --
    end process; 
    -- binary operator ADD_u2_u2_659_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_to_be_replaced_buffer, konst_658_wire_constant, tmp_var);
      ADD_u2_u2_659_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u2_u2_671_inst flow-through 
    process(ADD_u2_u2_671_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:ADD_u2_u2_671_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_670_wire_constant = "& Convert_SLV_To_Hex_String(konst_670_wire_constant) & " outputs:" & " ADD_u2_u2_671_wire= "  & Convert_SLV_To_Hex_String(ADD_u2_u2_671_wire));
      --
    end process; 
    -- binary operator ADD_u2_u2_671_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_to_be_replaced_buffer, konst_670_wire_constant, tmp_var);
      ADD_u2_u2_671_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_640_inst flow-through 
    process(EQ_u2_u1_640_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:EQ_u2_u1_640_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_639_wire_constant = "& Convert_SLV_To_Hex_String(konst_639_wire_constant) & " outputs:" & " EQ_u2_u1_640_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_640_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_640_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_to_be_replaced_buffer, konst_639_wire_constant, tmp_var);
      EQ_u2_u1_640_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_666_inst flow-through 
    process(EQ_u2_u1_666_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:EQ_u2_u1_666_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_665_wire_constant = "& Convert_SLV_To_Hex_String(konst_665_wire_constant) & " outputs:" & " EQ_u2_u1_666_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_666_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_666_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_to_be_replaced_buffer, konst_665_wire_constant, tmp_var);
      EQ_u2_u1_666_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_682_inst flow-through 
    process(MUL_u16_u16_682_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_682_inst:flowthrough inputs: " & " array_obj_ref_678_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_678_wire) & " array_obj_ref_681_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_681_wire) & " outputs:" & " MUL_u16_u16_682_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_682_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_682_inst
    process(array_obj_ref_678_wire, array_obj_ref_681_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_678_wire, array_obj_ref_681_wire, tmp_var);
      MUL_u16_u16_682_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_692_inst flow-through 
    process(MUL_u16_u16_692_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_692_inst:flowthrough inputs: " & " array_obj_ref_688_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_688_wire) & " array_obj_ref_691_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_691_wire) & " outputs:" & " MUL_u16_u16_692_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_692_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_692_inst
    process(array_obj_ref_688_wire, array_obj_ref_691_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_688_wire, array_obj_ref_691_wire, tmp_var);
      MUL_u16_u16_692_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_702_inst flow-through 
    process(MUL_u16_u16_702_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_702_inst:flowthrough inputs: " & " array_obj_ref_698_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_698_wire) & " array_obj_ref_701_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_701_wire) & " outputs:" & " MUL_u16_u16_702_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_702_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_702_inst
    process(array_obj_ref_698_wire, array_obj_ref_701_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_698_wire, array_obj_ref_701_wire, tmp_var);
      MUL_u16_u16_702_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_712_inst flow-through 
    process(MUL_u16_u16_712_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_712_inst:flowthrough inputs: " & " array_obj_ref_708_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_708_wire) & " array_obj_ref_711_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_711_wire) & " outputs:" & " MUL_u16_u16_712_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_712_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_712_inst
    process(array_obj_ref_708_wire, array_obj_ref_711_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_708_wire, array_obj_ref_711_wire, tmp_var);
      MUL_u16_u16_712_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_722_inst flow-through 
    process(MUL_u16_u16_722_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_722_inst:flowthrough inputs: " & " array_obj_ref_718_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_718_wire) & " array_obj_ref_721_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_721_wire) & " outputs:" & " MUL_u16_u16_722_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_722_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_722_inst
    process(array_obj_ref_718_wire, array_obj_ref_721_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_718_wire, array_obj_ref_721_wire, tmp_var);
      MUL_u16_u16_722_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_732_inst flow-through 
    process(MUL_u16_u16_732_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_732_inst:flowthrough inputs: " & " array_obj_ref_728_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_728_wire) & " array_obj_ref_731_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_731_wire) & " outputs:" & " MUL_u16_u16_732_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_732_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_732_inst
    process(array_obj_ref_728_wire, array_obj_ref_731_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_728_wire, array_obj_ref_731_wire, tmp_var);
      MUL_u16_u16_732_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_742_inst flow-through 
    process(MUL_u16_u16_742_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_742_inst:flowthrough inputs: " & " array_obj_ref_738_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_738_wire) & " array_obj_ref_741_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_741_wire) & " outputs:" & " MUL_u16_u16_742_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_742_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_742_inst
    process(array_obj_ref_738_wire, array_obj_ref_741_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_738_wire, array_obj_ref_741_wire, tmp_var);
      MUL_u16_u16_742_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_752_inst flow-through 
    process(MUL_u16_u16_752_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_752_inst:flowthrough inputs: " & " array_obj_ref_748_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_748_wire) & " array_obj_ref_751_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_751_wire) & " outputs:" & " MUL_u16_u16_752_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_752_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_752_inst
    process(array_obj_ref_748_wire, array_obj_ref_751_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_748_wire, array_obj_ref_751_wire, tmp_var);
      MUL_u16_u16_752_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_762_inst flow-through 
    process(MUL_u16_u16_762_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_762_inst:flowthrough inputs: " & " array_obj_ref_758_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_758_wire) & " array_obj_ref_761_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_761_wire) & " outputs:" & " MUL_u16_u16_762_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_762_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_762_inst
    process(array_obj_ref_758_wire, array_obj_ref_761_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_758_wire, array_obj_ref_761_wire, tmp_var);
      MUL_u16_u16_762_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_772_inst flow-through 
    process(MUL_u16_u16_772_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_772_inst:flowthrough inputs: " & " array_obj_ref_768_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_768_wire) & " array_obj_ref_771_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_771_wire) & " outputs:" & " MUL_u16_u16_772_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_772_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_772_inst
    process(array_obj_ref_768_wire, array_obj_ref_771_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_768_wire, array_obj_ref_771_wire, tmp_var);
      MUL_u16_u16_772_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_782_inst flow-through 
    process(MUL_u16_u16_782_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_782_inst:flowthrough inputs: " & " array_obj_ref_778_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_778_wire) & " array_obj_ref_781_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_781_wire) & " outputs:" & " MUL_u16_u16_782_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_782_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_782_inst
    process(array_obj_ref_778_wire, array_obj_ref_781_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_778_wire, array_obj_ref_781_wire, tmp_var);
      MUL_u16_u16_782_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_792_inst flow-through 
    process(MUL_u16_u16_792_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_792_inst:flowthrough inputs: " & " array_obj_ref_788_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_788_wire) & " array_obj_ref_791_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_791_wire) & " outputs:" & " MUL_u16_u16_792_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_792_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_792_inst
    process(array_obj_ref_788_wire, array_obj_ref_791_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_788_wire, array_obj_ref_791_wire, tmp_var);
      MUL_u16_u16_792_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_802_inst flow-through 
    process(MUL_u16_u16_802_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_802_inst:flowthrough inputs: " & " array_obj_ref_798_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_798_wire) & " array_obj_ref_801_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_801_wire) & " outputs:" & " MUL_u16_u16_802_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_802_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_802_inst
    process(array_obj_ref_798_wire, array_obj_ref_801_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_798_wire, array_obj_ref_801_wire, tmp_var);
      MUL_u16_u16_802_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_812_inst flow-through 
    process(MUL_u16_u16_812_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_812_inst:flowthrough inputs: " & " array_obj_ref_808_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_808_wire) & " array_obj_ref_811_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_811_wire) & " outputs:" & " MUL_u16_u16_812_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_812_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_812_inst
    process(array_obj_ref_808_wire, array_obj_ref_811_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_808_wire, array_obj_ref_811_wire, tmp_var);
      MUL_u16_u16_812_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_822_inst flow-through 
    process(MUL_u16_u16_822_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_822_inst:flowthrough inputs: " & " array_obj_ref_818_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_818_wire) & " array_obj_ref_821_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_821_wire) & " outputs:" & " MUL_u16_u16_822_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_822_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_822_inst
    process(array_obj_ref_818_wire, array_obj_ref_821_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_818_wire, array_obj_ref_821_wire, tmp_var);
      MUL_u16_u16_822_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_832_inst flow-through 
    process(MUL_u16_u16_832_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:MUL_u16_u16_832_inst:flowthrough inputs: " & " array_obj_ref_828_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_828_wire) & " array_obj_ref_831_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_831_wire) & " outputs:" & " MUL_u16_u16_832_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_832_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_832_inst
    process(array_obj_ref_828_wire, array_obj_ref_831_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_828_wire, array_obj_ref_831_wire, tmp_var);
      MUL_u16_u16_832_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u2_u2_645_inst flow-through 
    process(SUB_u2_u2_645_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:SUB_u2_u2_645_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_644_wire_constant = "& Convert_SLV_To_Hex_String(konst_644_wire_constant) & " outputs:" & " SUB_u2_u2_645_wire= "  & Convert_SLV_To_Hex_String(SUB_u2_u2_645_wire));
      --
    end process; 
    -- binary operator SUB_u2_u2_645_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntSub_proc(col_to_be_replaced_buffer, konst_644_wire_constant, tmp_var);
      SUB_u2_u2_645_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u2_u2_655_inst flow-through 
    process(SUB_u2_u2_655_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:SUB_u2_u2_655_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_654_wire_constant = "& Convert_SLV_To_Hex_String(konst_654_wire_constant) & " outputs:" & " SUB_u2_u2_655_wire= "  & Convert_SLV_To_Hex_String(SUB_u2_u2_655_wire));
      --
    end process; 
    -- binary operator SUB_u2_u2_655_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntSub_proc(col_to_be_replaced_buffer, konst_654_wire_constant, tmp_var);
      SUB_u2_u2_655_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGE_u2_u1_652_inst flow-through 
    process(UGE_u2_u1_652_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:UGE_u2_u1_652_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_651_wire_constant = "& Convert_SLV_To_Hex_String(konst_651_wire_constant) & " outputs:" & " UGE_u2_u1_652_wire= "  & Convert_SLV_To_Hex_String(UGE_u2_u1_652_wire));
      --
    end process; 
    -- binary operator UGE_u2_u1_652_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(col_to_be_replaced_buffer, konst_651_wire_constant, tmp_var);
      UGE_u2_u1_652_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_678_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_678_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_index_offset:started:   inputs: " & " R_col_to_be_replaced_677_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_677_scaled) & " array_obj_ref_678_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_678_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_678_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_index_offset:finished:  outputs: " & " array_obj_ref_678_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_678_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (38) : array_obj_ref_678_index_offset 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_677_scaled;
      array_obj_ref_678_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_678_index_offset_req_0;
      array_obj_ref_678_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_678_index_offset_req_1;
      array_obj_ref_678_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- logger for split-operator array_obj_ref_688_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_688_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_index_offset:started:   inputs: " & " R_col_to_be_replaced_687_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_687_scaled) & " array_obj_ref_688_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_688_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_688_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_index_offset:finished:  outputs: " & " array_obj_ref_688_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_688_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (39) : array_obj_ref_688_index_offset 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_687_scaled;
      array_obj_ref_688_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_688_index_offset_req_0;
      array_obj_ref_688_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_688_index_offset_req_1;
      array_obj_ref_688_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- logger for split-operator array_obj_ref_698_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_698_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_index_offset:started:   inputs: " & " R_col_to_be_replaced_697_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_697_scaled) & " array_obj_ref_698_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_698_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_698_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_index_offset:finished:  outputs: " & " array_obj_ref_698_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_698_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (40) : array_obj_ref_698_index_offset 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_697_scaled;
      array_obj_ref_698_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_698_index_offset_req_0;
      array_obj_ref_698_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_698_index_offset_req_1;
      array_obj_ref_698_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_40_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_40_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- logger for split-operator array_obj_ref_708_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_708_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_index_offset:started:   inputs: " & " R_col_to_be_replaced_707_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_707_scaled) & " array_obj_ref_708_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_708_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_708_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_index_offset:finished:  outputs: " & " array_obj_ref_708_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_708_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (41) : array_obj_ref_708_index_offset 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_707_scaled;
      array_obj_ref_708_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_708_index_offset_req_0;
      array_obj_ref_708_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_708_index_offset_req_1;
      array_obj_ref_708_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- logger for split-operator array_obj_ref_718_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_718_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_717_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_717_scaled) & " array_obj_ref_718_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_718_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_718_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_index_offset:finished:  outputs: " & " array_obj_ref_718_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_718_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (42) : array_obj_ref_718_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_717_scaled;
      array_obj_ref_718_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_718_index_offset_req_0;
      array_obj_ref_718_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_718_index_offset_req_1;
      array_obj_ref_718_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- logger for split-operator array_obj_ref_728_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_728_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_727_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_727_scaled) & " array_obj_ref_728_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_728_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_728_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_index_offset:finished:  outputs: " & " array_obj_ref_728_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_728_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (43) : array_obj_ref_728_index_offset 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_727_scaled;
      array_obj_ref_728_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_728_index_offset_req_0;
      array_obj_ref_728_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_728_index_offset_req_1;
      array_obj_ref_728_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- logger for split-operator array_obj_ref_738_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_738_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_737_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_737_scaled) & " array_obj_ref_738_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_738_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_738_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_index_offset:finished:  outputs: " & " array_obj_ref_738_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_738_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (44) : array_obj_ref_738_index_offset 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_737_scaled;
      array_obj_ref_738_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_738_index_offset_req_0;
      array_obj_ref_738_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_738_index_offset_req_1;
      array_obj_ref_738_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- logger for split-operator array_obj_ref_748_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_748_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_747_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_747_scaled) & " array_obj_ref_748_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_748_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_748_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_index_offset:finished:  outputs: " & " array_obj_ref_748_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_748_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (45) : array_obj_ref_748_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_747_scaled;
      array_obj_ref_748_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_748_index_offset_req_0;
      array_obj_ref_748_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_748_index_offset_req_1;
      array_obj_ref_748_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- logger for split-operator array_obj_ref_758_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_758_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_757_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_757_scaled) & " array_obj_ref_758_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_758_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_758_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_index_offset:finished:  outputs: " & " array_obj_ref_758_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_758_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (46) : array_obj_ref_758_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_757_scaled;
      array_obj_ref_758_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_758_index_offset_req_0;
      array_obj_ref_758_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_758_index_offset_req_1;
      array_obj_ref_758_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- logger for split-operator array_obj_ref_768_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_768_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_767_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_767_scaled) & " array_obj_ref_768_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_768_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_768_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_index_offset:finished:  outputs: " & " array_obj_ref_768_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_768_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (47) : array_obj_ref_768_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_767_scaled;
      array_obj_ref_768_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_768_index_offset_req_0;
      array_obj_ref_768_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_768_index_offset_req_1;
      array_obj_ref_768_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- logger for split-operator array_obj_ref_778_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_778_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_777_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_777_scaled) & " array_obj_ref_778_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_778_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_778_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_index_offset:finished:  outputs: " & " array_obj_ref_778_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_778_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (48) : array_obj_ref_778_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_777_scaled;
      array_obj_ref_778_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_778_index_offset_req_0;
      array_obj_ref_778_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_778_index_offset_req_1;
      array_obj_ref_778_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- logger for split-operator array_obj_ref_788_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_788_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_787_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_787_scaled) & " array_obj_ref_788_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_788_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_788_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_index_offset:finished:  outputs: " & " array_obj_ref_788_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_788_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (49) : array_obj_ref_788_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_787_scaled;
      array_obj_ref_788_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_788_index_offset_req_0;
      array_obj_ref_788_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_788_index_offset_req_1;
      array_obj_ref_788_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- logger for split-operator array_obj_ref_798_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_798_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_797_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_797_scaled) & " array_obj_ref_798_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_798_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_798_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_index_offset:finished:  outputs: " & " array_obj_ref_798_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_798_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (50) : array_obj_ref_798_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_797_scaled;
      array_obj_ref_798_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_798_index_offset_req_0;
      array_obj_ref_798_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_798_index_offset_req_1;
      array_obj_ref_798_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- logger for split-operator array_obj_ref_808_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_808_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_807_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_807_scaled) & " array_obj_ref_808_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_808_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_808_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_index_offset:finished:  outputs: " & " array_obj_ref_808_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_808_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (51) : array_obj_ref_808_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_807_scaled;
      array_obj_ref_808_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_808_index_offset_req_0;
      array_obj_ref_808_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_808_index_offset_req_1;
      array_obj_ref_808_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- logger for split-operator array_obj_ref_818_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_818_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_817_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_817_scaled) & " array_obj_ref_818_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_818_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_818_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_index_offset:finished:  outputs: " & " array_obj_ref_818_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_818_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (52) : array_obj_ref_818_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_817_scaled;
      array_obj_ref_818_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_818_index_offset_req_0;
      array_obj_ref_818_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_818_index_offset_req_1;
      array_obj_ref_818_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- logger for split-operator array_obj_ref_828_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_828_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_827_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_827_scaled) & " array_obj_ref_828_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_828_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_828_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_index_offset:finished:  outputs: " & " array_obj_ref_828_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_828_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (53) : array_obj_ref_828_index_offset 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_827_scaled;
      array_obj_ref_828_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_828_index_offset_req_0;
      array_obj_ref_828_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_828_index_offset_req_1;
      array_obj_ref_828_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- logger for split-operator array_obj_ref_688_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_688_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_load_0:started:   inputs: " & " array_obj_ref_688_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_688_word_address_0));
          --
        end if; 
        if array_obj_ref_688_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_688_load_0:finished:  outputs: " & " array_obj_ref_688_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_688_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_698_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_698_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_load_0:started:   inputs: " & " array_obj_ref_698_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_698_word_address_0));
          --
        end if; 
        if array_obj_ref_698_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_698_load_0:finished:  outputs: " & " array_obj_ref_698_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_698_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_738_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_738_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_load_0:started:   inputs: " & " array_obj_ref_738_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_738_word_address_0));
          --
        end if; 
        if array_obj_ref_738_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_738_load_0:finished:  outputs: " & " array_obj_ref_738_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_738_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_708_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_708_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_load_0:started:   inputs: " & " array_obj_ref_708_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_708_word_address_0));
          --
        end if; 
        if array_obj_ref_708_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_708_load_0:finished:  outputs: " & " array_obj_ref_708_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_708_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_678_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_678_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_load_0:started:   inputs: " & " array_obj_ref_678_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_678_word_address_0));
          --
        end if; 
        if array_obj_ref_678_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_678_load_0:finished:  outputs: " & " array_obj_ref_678_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_678_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_728_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_728_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_load_0:started:   inputs: " & " array_obj_ref_728_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_728_word_address_0));
          --
        end if; 
        if array_obj_ref_728_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_728_load_0:finished:  outputs: " & " array_obj_ref_728_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_728_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_718_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_718_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_load_0:started:   inputs: " & " array_obj_ref_718_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_718_word_address_0));
          --
        end if; 
        if array_obj_ref_718_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_718_load_0:finished:  outputs: " & " array_obj_ref_718_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_718_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_748_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_748_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_load_0:started:   inputs: " & " array_obj_ref_748_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_748_word_address_0));
          --
        end if; 
        if array_obj_ref_748_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_748_load_0:finished:  outputs: " & " array_obj_ref_748_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_748_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_758_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_758_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_load_0:started:   inputs: " & " array_obj_ref_758_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_758_word_address_0));
          --
        end if; 
        if array_obj_ref_758_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_758_load_0:finished:  outputs: " & " array_obj_ref_758_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_758_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_768_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_768_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_load_0:started:   inputs: " & " array_obj_ref_768_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_768_word_address_0));
          --
        end if; 
        if array_obj_ref_768_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_768_load_0:finished:  outputs: " & " array_obj_ref_768_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_768_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_778_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_778_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_load_0:started:   inputs: " & " array_obj_ref_778_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_778_word_address_0));
          --
        end if; 
        if array_obj_ref_778_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_778_load_0:finished:  outputs: " & " array_obj_ref_778_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_778_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_788_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_788_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_load_0:started:   inputs: " & " array_obj_ref_788_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_788_word_address_0));
          --
        end if; 
        if array_obj_ref_788_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_788_load_0:finished:  outputs: " & " array_obj_ref_788_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_788_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_798_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_798_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_load_0:started:   inputs: " & " array_obj_ref_798_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_798_word_address_0));
          --
        end if; 
        if array_obj_ref_798_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_798_load_0:finished:  outputs: " & " array_obj_ref_798_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_798_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_808_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_808_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_load_0:started:   inputs: " & " array_obj_ref_808_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_808_word_address_0));
          --
        end if; 
        if array_obj_ref_808_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_808_load_0:finished:  outputs: " & " array_obj_ref_808_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_808_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_818_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_818_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_load_0:started:   inputs: " & " array_obj_ref_818_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_818_word_address_0));
          --
        end if; 
        if array_obj_ref_818_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_818_load_0:finished:  outputs: " & " array_obj_ref_818_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_818_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_828_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_828_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_load_0:started:   inputs: " & " array_obj_ref_828_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_828_word_address_0));
          --
        end if; 
        if array_obj_ref_828_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_828_load_0:finished:  outputs: " & " array_obj_ref_828_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_828_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_688_load_0 array_obj_ref_698_load_0 array_obj_ref_738_load_0 array_obj_ref_708_load_0 array_obj_ref_678_load_0 array_obj_ref_728_load_0 array_obj_ref_718_load_0 array_obj_ref_748_load_0 array_obj_ref_758_load_0 array_obj_ref_768_load_0 array_obj_ref_778_load_0 array_obj_ref_788_load_0 array_obj_ref_798_load_0 array_obj_ref_808_load_0 array_obj_ref_818_load_0 array_obj_ref_828_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_688_load_0_req_0,
        array_obj_ref_688_load_0_ack_0,
        array_obj_ref_688_load_0_req_1,
        array_obj_ref_688_load_0_ack_1,
        "array_obj_ref_688_load_0",
        "memory_space_1" ,
        array_obj_ref_688_data_0,
        array_obj_ref_688_word_address_0,
        "array_obj_ref_688_data_0",
        "array_obj_ref_688_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_698_load_0_req_0,
        array_obj_ref_698_load_0_ack_0,
        array_obj_ref_698_load_0_req_1,
        array_obj_ref_698_load_0_ack_1,
        "array_obj_ref_698_load_0",
        "memory_space_1" ,
        array_obj_ref_698_data_0,
        array_obj_ref_698_word_address_0,
        "array_obj_ref_698_data_0",
        "array_obj_ref_698_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_738_load_0_req_0,
        array_obj_ref_738_load_0_ack_0,
        array_obj_ref_738_load_0_req_1,
        array_obj_ref_738_load_0_ack_1,
        "array_obj_ref_738_load_0",
        "memory_space_1" ,
        array_obj_ref_738_data_0,
        array_obj_ref_738_word_address_0,
        "array_obj_ref_738_data_0",
        "array_obj_ref_738_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_708_load_0_req_0,
        array_obj_ref_708_load_0_ack_0,
        array_obj_ref_708_load_0_req_1,
        array_obj_ref_708_load_0_ack_1,
        "array_obj_ref_708_load_0",
        "memory_space_1" ,
        array_obj_ref_708_data_0,
        array_obj_ref_708_word_address_0,
        "array_obj_ref_708_data_0",
        "array_obj_ref_708_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_678_load_0_req_0,
        array_obj_ref_678_load_0_ack_0,
        array_obj_ref_678_load_0_req_1,
        array_obj_ref_678_load_0_ack_1,
        "array_obj_ref_678_load_0",
        "memory_space_1" ,
        array_obj_ref_678_data_0,
        array_obj_ref_678_word_address_0,
        "array_obj_ref_678_data_0",
        "array_obj_ref_678_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_728_load_0_req_0,
        array_obj_ref_728_load_0_ack_0,
        array_obj_ref_728_load_0_req_1,
        array_obj_ref_728_load_0_ack_1,
        "array_obj_ref_728_load_0",
        "memory_space_1" ,
        array_obj_ref_728_data_0,
        array_obj_ref_728_word_address_0,
        "array_obj_ref_728_data_0",
        "array_obj_ref_728_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_718_load_0_req_0,
        array_obj_ref_718_load_0_ack_0,
        array_obj_ref_718_load_0_req_1,
        array_obj_ref_718_load_0_ack_1,
        "array_obj_ref_718_load_0",
        "memory_space_1" ,
        array_obj_ref_718_data_0,
        array_obj_ref_718_word_address_0,
        "array_obj_ref_718_data_0",
        "array_obj_ref_718_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_748_load_0_req_0,
        array_obj_ref_748_load_0_ack_0,
        array_obj_ref_748_load_0_req_1,
        array_obj_ref_748_load_0_ack_1,
        "array_obj_ref_748_load_0",
        "memory_space_1" ,
        array_obj_ref_748_data_0,
        array_obj_ref_748_word_address_0,
        "array_obj_ref_748_data_0",
        "array_obj_ref_748_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_758_load_0_req_0,
        array_obj_ref_758_load_0_ack_0,
        array_obj_ref_758_load_0_req_1,
        array_obj_ref_758_load_0_ack_1,
        "array_obj_ref_758_load_0",
        "memory_space_1" ,
        array_obj_ref_758_data_0,
        array_obj_ref_758_word_address_0,
        "array_obj_ref_758_data_0",
        "array_obj_ref_758_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_768_load_0_req_0,
        array_obj_ref_768_load_0_ack_0,
        array_obj_ref_768_load_0_req_1,
        array_obj_ref_768_load_0_ack_1,
        "array_obj_ref_768_load_0",
        "memory_space_1" ,
        array_obj_ref_768_data_0,
        array_obj_ref_768_word_address_0,
        "array_obj_ref_768_data_0",
        "array_obj_ref_768_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_778_load_0_req_0,
        array_obj_ref_778_load_0_ack_0,
        array_obj_ref_778_load_0_req_1,
        array_obj_ref_778_load_0_ack_1,
        "array_obj_ref_778_load_0",
        "memory_space_1" ,
        array_obj_ref_778_data_0,
        array_obj_ref_778_word_address_0,
        "array_obj_ref_778_data_0",
        "array_obj_ref_778_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_788_load_0_req_0,
        array_obj_ref_788_load_0_ack_0,
        array_obj_ref_788_load_0_req_1,
        array_obj_ref_788_load_0_ack_1,
        "array_obj_ref_788_load_0",
        "memory_space_1" ,
        array_obj_ref_788_data_0,
        array_obj_ref_788_word_address_0,
        "array_obj_ref_788_data_0",
        "array_obj_ref_788_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_798_load_0_req_0,
        array_obj_ref_798_load_0_ack_0,
        array_obj_ref_798_load_0_req_1,
        array_obj_ref_798_load_0_ack_1,
        "array_obj_ref_798_load_0",
        "memory_space_1" ,
        array_obj_ref_798_data_0,
        array_obj_ref_798_word_address_0,
        "array_obj_ref_798_data_0",
        "array_obj_ref_798_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_808_load_0_req_0,
        array_obj_ref_808_load_0_ack_0,
        array_obj_ref_808_load_0_req_1,
        array_obj_ref_808_load_0_ack_1,
        "array_obj_ref_808_load_0",
        "memory_space_1" ,
        array_obj_ref_808_data_0,
        array_obj_ref_808_word_address_0,
        "array_obj_ref_808_data_0",
        "array_obj_ref_808_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_818_load_0_req_0,
        array_obj_ref_818_load_0_ack_0,
        array_obj_ref_818_load_0_req_1,
        array_obj_ref_818_load_0_ack_1,
        "array_obj_ref_818_load_0",
        "memory_space_1" ,
        array_obj_ref_818_data_0,
        array_obj_ref_818_word_address_0,
        "array_obj_ref_818_data_0",
        "array_obj_ref_818_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_828_load_0_req_0,
        array_obj_ref_828_load_0_ack_0,
        array_obj_ref_828_load_0_req_1,
        array_obj_ref_828_load_0_ack_1,
        "array_obj_ref_828_load_0",
        "memory_space_1" ,
        array_obj_ref_828_data_0,
        array_obj_ref_828_word_address_0,
        "array_obj_ref_828_data_0",
        "array_obj_ref_828_word_address_0" -- 
      );
      reqL_unguarded(15) <= array_obj_ref_688_load_0_req_0;
      reqL_unguarded(14) <= array_obj_ref_698_load_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_738_load_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_708_load_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_678_load_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_728_load_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_718_load_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_748_load_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_758_load_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_768_load_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_778_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_788_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_798_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_808_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_818_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_828_load_0_req_0;
      array_obj_ref_688_load_0_ack_0 <= ackL_unguarded(15);
      array_obj_ref_698_load_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_738_load_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_708_load_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_678_load_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_728_load_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_718_load_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_748_load_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_758_load_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_768_load_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_778_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_788_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_798_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_808_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_818_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_828_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= array_obj_ref_688_load_0_req_1;
      reqR_unguarded(14) <= array_obj_ref_698_load_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_738_load_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_708_load_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_678_load_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_728_load_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_718_load_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_748_load_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_758_load_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_768_load_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_778_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_788_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_798_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_808_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_818_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_828_load_0_req_1;
      array_obj_ref_688_load_0_ack_1 <= ackR_unguarded(15);
      array_obj_ref_698_load_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_738_load_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_708_load_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_678_load_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_728_load_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_718_load_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_748_load_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_758_load_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_768_load_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_778_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_788_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_798_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_808_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_818_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_828_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_688_word_address_0 & array_obj_ref_698_word_address_0 & array_obj_ref_738_word_address_0 & array_obj_ref_708_word_address_0 & array_obj_ref_678_word_address_0 & array_obj_ref_728_word_address_0 & array_obj_ref_718_word_address_0 & array_obj_ref_748_word_address_0 & array_obj_ref_758_word_address_0 & array_obj_ref_768_word_address_0 & array_obj_ref_778_word_address_0 & array_obj_ref_788_word_address_0 & array_obj_ref_798_word_address_0 & array_obj_ref_808_word_address_0 & array_obj_ref_818_word_address_0 & array_obj_ref_828_word_address_0;
      array_obj_ref_688_data_0 <= data_out(255 downto 240);
      array_obj_ref_698_data_0 <= data_out(239 downto 224);
      array_obj_ref_738_data_0 <= data_out(223 downto 208);
      array_obj_ref_708_data_0 <= data_out(207 downto 192);
      array_obj_ref_678_data_0 <= data_out(191 downto 176);
      array_obj_ref_728_data_0 <= data_out(175 downto 160);
      array_obj_ref_718_data_0 <= data_out(159 downto 144);
      array_obj_ref_748_data_0 <= data_out(143 downto 128);
      array_obj_ref_758_data_0 <= data_out(127 downto 112);
      array_obj_ref_768_data_0 <= data_out(111 downto 96);
      array_obj_ref_778_data_0 <= data_out(95 downto 80);
      array_obj_ref_788_data_0 <= data_out(79 downto 64);
      array_obj_ref_798_data_0 <= data_out(63 downto 48);
      array_obj_ref_808_data_0 <= data_out(47 downto 32);
      array_obj_ref_818_data_0 <= data_out(31 downto 16);
      array_obj_ref_828_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 4,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(3 downto 0),
          mtag => memory_space_1_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_701_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_701_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_701_load_0:started:   inputs: " & " array_obj_ref_701_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_701_word_address_0));
          --
        end if; 
        if array_obj_ref_701_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_701_load_0:finished:  outputs: " & " array_obj_ref_701_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_701_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_691_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_691_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_691_load_0:started:   inputs: " & " array_obj_ref_691_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_691_word_address_0));
          --
        end if; 
        if array_obj_ref_691_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_691_load_0:finished:  outputs: " & " array_obj_ref_691_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_691_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_711_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_711_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_711_load_0:started:   inputs: " & " array_obj_ref_711_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_711_word_address_0));
          --
        end if; 
        if array_obj_ref_711_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_711_load_0:finished:  outputs: " & " array_obj_ref_711_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_711_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_681_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_681_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_681_load_0:started:   inputs: " & " array_obj_ref_681_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_681_word_address_0));
          --
        end if; 
        if array_obj_ref_681_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_681_load_0:finished:  outputs: " & " array_obj_ref_681_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_681_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_731_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_731_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_731_load_0:started:   inputs: " & " array_obj_ref_731_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_731_word_address_0));
          --
        end if; 
        if array_obj_ref_731_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_731_load_0:finished:  outputs: " & " array_obj_ref_731_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_731_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_721_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_721_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_721_load_0:started:   inputs: " & " array_obj_ref_721_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_721_word_address_0));
          --
        end if; 
        if array_obj_ref_721_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_721_load_0:finished:  outputs: " & " array_obj_ref_721_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_721_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_741_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_741_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_741_load_0:started:   inputs: " & " array_obj_ref_741_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_741_word_address_0));
          --
        end if; 
        if array_obj_ref_741_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_741_load_0:finished:  outputs: " & " array_obj_ref_741_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_741_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_751_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_751_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_751_load_0:started:   inputs: " & " array_obj_ref_751_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_751_word_address_0));
          --
        end if; 
        if array_obj_ref_751_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_751_load_0:finished:  outputs: " & " array_obj_ref_751_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_751_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_761_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_761_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_761_load_0:started:   inputs: " & " array_obj_ref_761_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_761_word_address_0));
          --
        end if; 
        if array_obj_ref_761_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_761_load_0:finished:  outputs: " & " array_obj_ref_761_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_761_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_771_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_771_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_771_load_0:started:   inputs: " & " array_obj_ref_771_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_771_word_address_0));
          --
        end if; 
        if array_obj_ref_771_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_771_load_0:finished:  outputs: " & " array_obj_ref_771_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_771_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_781_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_781_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_781_load_0:started:   inputs: " & " array_obj_ref_781_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_781_word_address_0));
          --
        end if; 
        if array_obj_ref_781_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_781_load_0:finished:  outputs: " & " array_obj_ref_781_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_781_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_791_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_791_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_791_load_0:started:   inputs: " & " array_obj_ref_791_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_791_word_address_0));
          --
        end if; 
        if array_obj_ref_791_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_791_load_0:finished:  outputs: " & " array_obj_ref_791_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_791_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_801_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_801_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_801_load_0:started:   inputs: " & " array_obj_ref_801_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_801_word_address_0));
          --
        end if; 
        if array_obj_ref_801_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_801_load_0:finished:  outputs: " & " array_obj_ref_801_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_801_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_811_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_811_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_811_load_0:started:   inputs: " & " array_obj_ref_811_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_811_word_address_0));
          --
        end if; 
        if array_obj_ref_811_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_811_load_0:finished:  outputs: " & " array_obj_ref_811_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_811_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_821_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_821_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_821_load_0:started:   inputs: " & " array_obj_ref_821_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_821_word_address_0));
          --
        end if; 
        if array_obj_ref_821_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_821_load_0:finished:  outputs: " & " array_obj_ref_821_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_821_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_831_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_831_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_831_load_0:started:   inputs: " & " array_obj_ref_831_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_831_word_address_0));
          --
        end if; 
        if array_obj_ref_831_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc:DP:array_obj_ref_831_load_0:finished:  outputs: " & " array_obj_ref_831_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_831_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (1) : array_obj_ref_701_load_0 array_obj_ref_691_load_0 array_obj_ref_711_load_0 array_obj_ref_681_load_0 array_obj_ref_731_load_0 array_obj_ref_721_load_0 array_obj_ref_741_load_0 array_obj_ref_751_load_0 array_obj_ref_761_load_0 array_obj_ref_771_load_0 array_obj_ref_781_load_0 array_obj_ref_791_load_0 array_obj_ref_801_load_0 array_obj_ref_811_load_0 array_obj_ref_821_load_0 array_obj_ref_831_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_701_load_0_req_0,
        array_obj_ref_701_load_0_ack_0,
        array_obj_ref_701_load_0_req_1,
        array_obj_ref_701_load_0_ack_1,
        "array_obj_ref_701_load_0",
        "memory_space_0" ,
        array_obj_ref_701_data_0,
        array_obj_ref_701_word_address_0,
        "array_obj_ref_701_data_0",
        "array_obj_ref_701_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_691_load_0_req_0,
        array_obj_ref_691_load_0_ack_0,
        array_obj_ref_691_load_0_req_1,
        array_obj_ref_691_load_0_ack_1,
        "array_obj_ref_691_load_0",
        "memory_space_0" ,
        array_obj_ref_691_data_0,
        array_obj_ref_691_word_address_0,
        "array_obj_ref_691_data_0",
        "array_obj_ref_691_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_711_load_0_req_0,
        array_obj_ref_711_load_0_ack_0,
        array_obj_ref_711_load_0_req_1,
        array_obj_ref_711_load_0_ack_1,
        "array_obj_ref_711_load_0",
        "memory_space_0" ,
        array_obj_ref_711_data_0,
        array_obj_ref_711_word_address_0,
        "array_obj_ref_711_data_0",
        "array_obj_ref_711_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_681_load_0_req_0,
        array_obj_ref_681_load_0_ack_0,
        array_obj_ref_681_load_0_req_1,
        array_obj_ref_681_load_0_ack_1,
        "array_obj_ref_681_load_0",
        "memory_space_0" ,
        array_obj_ref_681_data_0,
        array_obj_ref_681_word_address_0,
        "array_obj_ref_681_data_0",
        "array_obj_ref_681_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_731_load_0_req_0,
        array_obj_ref_731_load_0_ack_0,
        array_obj_ref_731_load_0_req_1,
        array_obj_ref_731_load_0_ack_1,
        "array_obj_ref_731_load_0",
        "memory_space_0" ,
        array_obj_ref_731_data_0,
        array_obj_ref_731_word_address_0,
        "array_obj_ref_731_data_0",
        "array_obj_ref_731_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_721_load_0_req_0,
        array_obj_ref_721_load_0_ack_0,
        array_obj_ref_721_load_0_req_1,
        array_obj_ref_721_load_0_ack_1,
        "array_obj_ref_721_load_0",
        "memory_space_0" ,
        array_obj_ref_721_data_0,
        array_obj_ref_721_word_address_0,
        "array_obj_ref_721_data_0",
        "array_obj_ref_721_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_741_load_0_req_0,
        array_obj_ref_741_load_0_ack_0,
        array_obj_ref_741_load_0_req_1,
        array_obj_ref_741_load_0_ack_1,
        "array_obj_ref_741_load_0",
        "memory_space_0" ,
        array_obj_ref_741_data_0,
        array_obj_ref_741_word_address_0,
        "array_obj_ref_741_data_0",
        "array_obj_ref_741_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_751_load_0_req_0,
        array_obj_ref_751_load_0_ack_0,
        array_obj_ref_751_load_0_req_1,
        array_obj_ref_751_load_0_ack_1,
        "array_obj_ref_751_load_0",
        "memory_space_0" ,
        array_obj_ref_751_data_0,
        array_obj_ref_751_word_address_0,
        "array_obj_ref_751_data_0",
        "array_obj_ref_751_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_761_load_0_req_0,
        array_obj_ref_761_load_0_ack_0,
        array_obj_ref_761_load_0_req_1,
        array_obj_ref_761_load_0_ack_1,
        "array_obj_ref_761_load_0",
        "memory_space_0" ,
        array_obj_ref_761_data_0,
        array_obj_ref_761_word_address_0,
        "array_obj_ref_761_data_0",
        "array_obj_ref_761_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_771_load_0_req_0,
        array_obj_ref_771_load_0_ack_0,
        array_obj_ref_771_load_0_req_1,
        array_obj_ref_771_load_0_ack_1,
        "array_obj_ref_771_load_0",
        "memory_space_0" ,
        array_obj_ref_771_data_0,
        array_obj_ref_771_word_address_0,
        "array_obj_ref_771_data_0",
        "array_obj_ref_771_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_781_load_0_req_0,
        array_obj_ref_781_load_0_ack_0,
        array_obj_ref_781_load_0_req_1,
        array_obj_ref_781_load_0_ack_1,
        "array_obj_ref_781_load_0",
        "memory_space_0" ,
        array_obj_ref_781_data_0,
        array_obj_ref_781_word_address_0,
        "array_obj_ref_781_data_0",
        "array_obj_ref_781_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_791_load_0_req_0,
        array_obj_ref_791_load_0_ack_0,
        array_obj_ref_791_load_0_req_1,
        array_obj_ref_791_load_0_ack_1,
        "array_obj_ref_791_load_0",
        "memory_space_0" ,
        array_obj_ref_791_data_0,
        array_obj_ref_791_word_address_0,
        "array_obj_ref_791_data_0",
        "array_obj_ref_791_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_801_load_0_req_0,
        array_obj_ref_801_load_0_ack_0,
        array_obj_ref_801_load_0_req_1,
        array_obj_ref_801_load_0_ack_1,
        "array_obj_ref_801_load_0",
        "memory_space_0" ,
        array_obj_ref_801_data_0,
        array_obj_ref_801_word_address_0,
        "array_obj_ref_801_data_0",
        "array_obj_ref_801_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_811_load_0_req_0,
        array_obj_ref_811_load_0_ack_0,
        array_obj_ref_811_load_0_req_1,
        array_obj_ref_811_load_0_ack_1,
        "array_obj_ref_811_load_0",
        "memory_space_0" ,
        array_obj_ref_811_data_0,
        array_obj_ref_811_word_address_0,
        "array_obj_ref_811_data_0",
        "array_obj_ref_811_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_821_load_0_req_0,
        array_obj_ref_821_load_0_ack_0,
        array_obj_ref_821_load_0_req_1,
        array_obj_ref_821_load_0_ack_1,
        "array_obj_ref_821_load_0",
        "memory_space_0" ,
        array_obj_ref_821_data_0,
        array_obj_ref_821_word_address_0,
        "array_obj_ref_821_data_0",
        "array_obj_ref_821_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_831_load_0_req_0,
        array_obj_ref_831_load_0_ack_0,
        array_obj_ref_831_load_0_req_1,
        array_obj_ref_831_load_0_ack_1,
        "array_obj_ref_831_load_0",
        "memory_space_0" ,
        array_obj_ref_831_data_0,
        array_obj_ref_831_word_address_0,
        "array_obj_ref_831_data_0",
        "array_obj_ref_831_word_address_0" -- 
      );
      reqL_unguarded(15) <= array_obj_ref_701_load_0_req_0;
      reqL_unguarded(14) <= array_obj_ref_691_load_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_711_load_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_681_load_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_731_load_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_721_load_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_741_load_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_751_load_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_761_load_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_771_load_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_781_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_791_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_801_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_811_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_821_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_831_load_0_req_0;
      array_obj_ref_701_load_0_ack_0 <= ackL_unguarded(15);
      array_obj_ref_691_load_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_711_load_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_681_load_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_731_load_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_721_load_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_741_load_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_751_load_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_761_load_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_771_load_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_781_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_791_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_801_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_811_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_821_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_831_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= array_obj_ref_701_load_0_req_1;
      reqR_unguarded(14) <= array_obj_ref_691_load_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_711_load_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_681_load_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_731_load_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_721_load_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_741_load_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_751_load_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_761_load_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_771_load_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_781_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_791_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_801_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_811_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_821_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_831_load_0_req_1;
      array_obj_ref_701_load_0_ack_1 <= ackR_unguarded(15);
      array_obj_ref_691_load_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_711_load_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_681_load_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_731_load_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_721_load_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_741_load_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_751_load_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_761_load_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_771_load_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_781_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_791_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_801_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_811_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_821_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_831_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_701_word_address_0 & array_obj_ref_691_word_address_0 & array_obj_ref_711_word_address_0 & array_obj_ref_681_word_address_0 & array_obj_ref_731_word_address_0 & array_obj_ref_721_word_address_0 & array_obj_ref_741_word_address_0 & array_obj_ref_751_word_address_0 & array_obj_ref_761_word_address_0 & array_obj_ref_771_word_address_0 & array_obj_ref_781_word_address_0 & array_obj_ref_791_word_address_0 & array_obj_ref_801_word_address_0 & array_obj_ref_811_word_address_0 & array_obj_ref_821_word_address_0 & array_obj_ref_831_word_address_0;
      array_obj_ref_701_data_0 <= data_out(255 downto 240);
      array_obj_ref_691_data_0 <= data_out(239 downto 224);
      array_obj_ref_711_data_0 <= data_out(223 downto 208);
      array_obj_ref_681_data_0 <= data_out(207 downto 192);
      array_obj_ref_731_data_0 <= data_out(191 downto 176);
      array_obj_ref_721_data_0 <= data_out(175 downto 160);
      array_obj_ref_741_data_0 <= data_out(159 downto 144);
      array_obj_ref_751_data_0 <= data_out(143 downto 128);
      array_obj_ref_761_data_0 <= data_out(127 downto 112);
      array_obj_ref_771_data_0 <= data_out(111 downto 96);
      array_obj_ref_781_data_0 <= data_out(95 downto 80);
      array_obj_ref_791_data_0 <= data_out(79 downto 64);
      array_obj_ref_801_data_0 <= data_out(63 downto 48);
      array_obj_ref_811_data_0 <= data_out(47 downto 32);
      array_obj_ref_821_data_0 <= data_out(31 downto 16);
      array_obj_ref_831_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 4,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(3 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- 
  end Block; -- data_path
  -- 
end mainAcc_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity mainAcc2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    I : in  std_logic_vector(5 downto 0);
    J : in  std_logic_vector(4 downto 0);
    col_to_be_replaced : in  std_logic_vector(1 downto 0);
    ofmap_pixel : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mainAcc2;
architecture mainAcc2_arch of mainAcc2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 13)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal I_buffer :  std_logic_vector(5 downto 0);
  signal I_update_enable: Boolean;
  signal J_buffer :  std_logic_vector(4 downto 0);
  signal J_update_enable: Boolean;
  signal col_to_be_replaced_buffer :  std_logic_vector(1 downto 0);
  signal col_to_be_replaced_update_enable: Boolean;
  -- output port buffer signals
  signal ofmap_pixel_buffer :  std_logic_vector(15 downto 0);
  signal ofmap_pixel_update_enable: Boolean;
  signal mainAcc2_CP_4584_start: Boolean;
  signal mainAcc2_CP_4584_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1003_inst_ack_1 : boolean;
  signal array_obj_ref_998_index_offset_ack_0 : boolean;
  signal array_obj_ref_1008_load_0_req_1 : boolean;
  signal array_obj_ref_998_load_0_req_0 : boolean;
  signal type_cast_1003_inst_req_1 : boolean;
  signal array_obj_ref_1001_load_0_req_0 : boolean;
  signal array_obj_ref_1008_index_offset_req_1 : boolean;
  signal array_obj_ref_1098_load_0_req_0 : boolean;
  signal type_cast_993_inst_req_0 : boolean;
  signal array_obj_ref_1008_load_0_ack_0 : boolean;
  signal array_obj_ref_1008_load_0_req_0 : boolean;
  signal array_obj_ref_991_load_0_req_0 : boolean;
  signal array_obj_ref_988_index_offset_req_0 : boolean;
  signal type_cast_1003_inst_req_0 : boolean;
  signal type_cast_1003_inst_ack_0 : boolean;
  signal array_obj_ref_1008_index_offset_ack_1 : boolean;
  signal array_obj_ref_988_index_offset_ack_0 : boolean;
  signal array_obj_ref_988_index_offset_req_1 : boolean;
  signal array_obj_ref_998_load_0_req_1 : boolean;
  signal array_obj_ref_988_index_offset_ack_1 : boolean;
  signal array_obj_ref_998_load_0_ack_1 : boolean;
  signal array_obj_ref_988_load_0_req_0 : boolean;
  signal array_obj_ref_1008_load_0_ack_1 : boolean;
  signal array_obj_ref_988_load_0_req_1 : boolean;
  signal array_obj_ref_1098_load_0_ack_0 : boolean;
  signal array_obj_ref_988_load_0_ack_0 : boolean;
  signal array_obj_ref_988_load_0_ack_1 : boolean;
  signal array_obj_ref_991_load_0_req_1 : boolean;
  signal type_cast_993_inst_ack_0 : boolean;
  signal array_obj_ref_998_load_0_ack_0 : boolean;
  signal array_obj_ref_991_load_0_ack_1 : boolean;
  signal array_obj_ref_991_load_0_ack_0 : boolean;
  signal type_cast_993_inst_req_1 : boolean;
  signal array_obj_ref_998_index_offset_req_0 : boolean;
  signal array_obj_ref_1001_load_0_ack_0 : boolean;
  signal type_cast_993_inst_ack_1 : boolean;
  signal array_obj_ref_1011_load_0_req_0 : boolean;
  signal type_cast_1013_inst_req_1 : boolean;
  signal type_cast_1013_inst_ack_1 : boolean;
  signal type_cast_1013_inst_ack_0 : boolean;
  signal type_cast_1013_inst_req_0 : boolean;
  signal type_cast_1103_inst_req_1 : boolean;
  signal array_obj_ref_1011_load_0_req_1 : boolean;
  signal array_obj_ref_1011_load_0_ack_1 : boolean;
  signal type_cast_1103_inst_ack_1 : boolean;
  signal array_obj_ref_1011_load_0_ack_0 : boolean;
  signal array_obj_ref_1008_index_offset_ack_0 : boolean;
  signal array_obj_ref_1001_load_0_ack_1 : boolean;
  signal array_obj_ref_1008_index_offset_req_0 : boolean;
  signal array_obj_ref_998_index_offset_ack_1 : boolean;
  signal array_obj_ref_1001_load_0_req_1 : boolean;
  signal array_obj_ref_998_index_offset_req_1 : boolean;
  signal array_obj_ref_1108_index_offset_req_1 : boolean;
  signal array_obj_ref_1108_index_offset_ack_1 : boolean;
  signal MUX_957_inst_req_0 : boolean;
  signal MUX_957_inst_ack_0 : boolean;
  signal MUX_957_inst_req_1 : boolean;
  signal MUX_957_inst_ack_1 : boolean;
  signal MUX_971_inst_req_0 : boolean;
  signal MUX_971_inst_ack_0 : boolean;
  signal MUX_971_inst_req_1 : boolean;
  signal MUX_971_inst_ack_1 : boolean;
  signal MUX_983_inst_req_0 : boolean;
  signal MUX_983_inst_ack_0 : boolean;
  signal MUX_983_inst_req_1 : boolean;
  signal MUX_983_inst_ack_1 : boolean;
  signal array_obj_ref_1018_index_offset_req_0 : boolean;
  signal array_obj_ref_1018_index_offset_ack_0 : boolean;
  signal array_obj_ref_1018_index_offset_req_1 : boolean;
  signal array_obj_ref_1018_index_offset_ack_1 : boolean;
  signal array_obj_ref_1018_load_0_req_0 : boolean;
  signal array_obj_ref_1018_load_0_ack_0 : boolean;
  signal array_obj_ref_1018_load_0_req_1 : boolean;
  signal array_obj_ref_1018_load_0_ack_1 : boolean;
  signal array_obj_ref_1021_load_0_req_0 : boolean;
  signal array_obj_ref_1021_load_0_ack_0 : boolean;
  signal array_obj_ref_1021_load_0_req_1 : boolean;
  signal array_obj_ref_1021_load_0_ack_1 : boolean;
  signal type_cast_1023_inst_req_0 : boolean;
  signal type_cast_1023_inst_ack_0 : boolean;
  signal type_cast_1023_inst_req_1 : boolean;
  signal type_cast_1023_inst_ack_1 : boolean;
  signal array_obj_ref_1028_index_offset_req_0 : boolean;
  signal array_obj_ref_1028_index_offset_ack_0 : boolean;
  signal array_obj_ref_1028_index_offset_req_1 : boolean;
  signal array_obj_ref_1028_index_offset_ack_1 : boolean;
  signal array_obj_ref_1028_load_0_req_0 : boolean;
  signal array_obj_ref_1028_load_0_ack_0 : boolean;
  signal array_obj_ref_1028_load_0_req_1 : boolean;
  signal array_obj_ref_1028_load_0_ack_1 : boolean;
  signal array_obj_ref_1031_load_0_req_0 : boolean;
  signal array_obj_ref_1031_load_0_ack_0 : boolean;
  signal array_obj_ref_1031_load_0_req_1 : boolean;
  signal array_obj_ref_1031_load_0_ack_1 : boolean;
  signal type_cast_1033_inst_req_0 : boolean;
  signal type_cast_1033_inst_ack_0 : boolean;
  signal type_cast_1033_inst_req_1 : boolean;
  signal type_cast_1033_inst_ack_1 : boolean;
  signal array_obj_ref_1038_index_offset_req_0 : boolean;
  signal array_obj_ref_1038_index_offset_ack_0 : boolean;
  signal array_obj_ref_1038_index_offset_req_1 : boolean;
  signal array_obj_ref_1038_index_offset_ack_1 : boolean;
  signal array_obj_ref_1038_load_0_req_0 : boolean;
  signal array_obj_ref_1038_load_0_ack_0 : boolean;
  signal array_obj_ref_1038_load_0_req_1 : boolean;
  signal array_obj_ref_1038_load_0_ack_1 : boolean;
  signal array_obj_ref_1041_load_0_req_0 : boolean;
  signal array_obj_ref_1041_load_0_ack_0 : boolean;
  signal array_obj_ref_1041_load_0_req_1 : boolean;
  signal array_obj_ref_1041_load_0_ack_1 : boolean;
  signal type_cast_1043_inst_req_0 : boolean;
  signal type_cast_1043_inst_ack_0 : boolean;
  signal type_cast_1043_inst_req_1 : boolean;
  signal type_cast_1043_inst_ack_1 : boolean;
  signal type_cast_1103_inst_ack_0 : boolean;
  signal array_obj_ref_1048_index_offset_req_0 : boolean;
  signal array_obj_ref_1048_index_offset_ack_0 : boolean;
  signal type_cast_1103_inst_req_0 : boolean;
  signal array_obj_ref_1048_index_offset_req_1 : boolean;
  signal array_obj_ref_1048_index_offset_ack_1 : boolean;
  signal array_obj_ref_1048_load_0_req_0 : boolean;
  signal array_obj_ref_1048_load_0_ack_0 : boolean;
  signal array_obj_ref_1101_load_0_ack_1 : boolean;
  signal array_obj_ref_1101_load_0_req_1 : boolean;
  signal array_obj_ref_1048_load_0_req_1 : boolean;
  signal array_obj_ref_1048_load_0_ack_1 : boolean;
  signal array_obj_ref_1108_index_offset_req_0 : boolean;
  signal array_obj_ref_1108_index_offset_ack_0 : boolean;
  signal array_obj_ref_1051_load_0_req_0 : boolean;
  signal array_obj_ref_1051_load_0_ack_0 : boolean;
  signal array_obj_ref_1101_load_0_ack_0 : boolean;
  signal array_obj_ref_1051_load_0_req_1 : boolean;
  signal array_obj_ref_1051_load_0_ack_1 : boolean;
  signal array_obj_ref_1101_load_0_req_0 : boolean;
  signal type_cast_1053_inst_req_0 : boolean;
  signal type_cast_1053_inst_ack_0 : boolean;
  signal type_cast_1053_inst_req_1 : boolean;
  signal type_cast_1053_inst_ack_1 : boolean;
  signal array_obj_ref_1058_index_offset_req_0 : boolean;
  signal array_obj_ref_1058_index_offset_ack_0 : boolean;
  signal array_obj_ref_1058_index_offset_req_1 : boolean;
  signal array_obj_ref_1058_index_offset_ack_1 : boolean;
  signal array_obj_ref_1058_load_0_req_0 : boolean;
  signal array_obj_ref_1058_load_0_ack_0 : boolean;
  signal array_obj_ref_1058_load_0_req_1 : boolean;
  signal array_obj_ref_1058_load_0_ack_1 : boolean;
  signal array_obj_ref_1098_load_0_ack_1 : boolean;
  signal array_obj_ref_1061_load_0_req_0 : boolean;
  signal array_obj_ref_1061_load_0_ack_0 : boolean;
  signal array_obj_ref_1098_load_0_req_1 : boolean;
  signal array_obj_ref_1061_load_0_req_1 : boolean;
  signal array_obj_ref_1061_load_0_ack_1 : boolean;
  signal type_cast_1063_inst_req_0 : boolean;
  signal type_cast_1063_inst_ack_0 : boolean;
  signal type_cast_1063_inst_req_1 : boolean;
  signal type_cast_1063_inst_ack_1 : boolean;
  signal array_obj_ref_1068_index_offset_req_0 : boolean;
  signal array_obj_ref_1068_index_offset_ack_0 : boolean;
  signal array_obj_ref_1068_index_offset_req_1 : boolean;
  signal array_obj_ref_1068_index_offset_ack_1 : boolean;
  signal array_obj_ref_1068_load_0_req_0 : boolean;
  signal array_obj_ref_1068_load_0_ack_0 : boolean;
  signal array_obj_ref_1068_load_0_req_1 : boolean;
  signal array_obj_ref_1068_load_0_ack_1 : boolean;
  signal array_obj_ref_1071_load_0_req_0 : boolean;
  signal array_obj_ref_1071_load_0_ack_0 : boolean;
  signal array_obj_ref_1071_load_0_req_1 : boolean;
  signal array_obj_ref_1071_load_0_ack_1 : boolean;
  signal type_cast_1073_inst_req_0 : boolean;
  signal type_cast_1073_inst_ack_0 : boolean;
  signal type_cast_1073_inst_req_1 : boolean;
  signal type_cast_1073_inst_ack_1 : boolean;
  signal array_obj_ref_1078_index_offset_req_0 : boolean;
  signal array_obj_ref_1078_index_offset_ack_0 : boolean;
  signal array_obj_ref_1078_index_offset_req_1 : boolean;
  signal array_obj_ref_1078_index_offset_ack_1 : boolean;
  signal array_obj_ref_1078_load_0_req_0 : boolean;
  signal array_obj_ref_1078_load_0_ack_0 : boolean;
  signal array_obj_ref_1078_load_0_req_1 : boolean;
  signal array_obj_ref_1078_load_0_ack_1 : boolean;
  signal array_obj_ref_1081_load_0_req_0 : boolean;
  signal array_obj_ref_1081_load_0_ack_0 : boolean;
  signal array_obj_ref_1081_load_0_req_1 : boolean;
  signal array_obj_ref_1081_load_0_ack_1 : boolean;
  signal type_cast_1083_inst_req_0 : boolean;
  signal type_cast_1083_inst_ack_0 : boolean;
  signal type_cast_1083_inst_req_1 : boolean;
  signal type_cast_1083_inst_ack_1 : boolean;
  signal array_obj_ref_1088_index_offset_req_0 : boolean;
  signal array_obj_ref_1088_index_offset_ack_0 : boolean;
  signal array_obj_ref_1088_index_offset_req_1 : boolean;
  signal array_obj_ref_1088_index_offset_ack_1 : boolean;
  signal array_obj_ref_1088_load_0_req_0 : boolean;
  signal array_obj_ref_1088_load_0_ack_0 : boolean;
  signal array_obj_ref_1088_load_0_req_1 : boolean;
  signal array_obj_ref_1088_load_0_ack_1 : boolean;
  signal array_obj_ref_1091_load_0_req_0 : boolean;
  signal array_obj_ref_1091_load_0_ack_0 : boolean;
  signal array_obj_ref_1091_load_0_req_1 : boolean;
  signal array_obj_ref_1091_load_0_ack_1 : boolean;
  signal type_cast_1093_inst_req_0 : boolean;
  signal type_cast_1093_inst_ack_0 : boolean;
  signal type_cast_1093_inst_req_1 : boolean;
  signal type_cast_1093_inst_ack_1 : boolean;
  signal array_obj_ref_1098_index_offset_req_0 : boolean;
  signal array_obj_ref_1098_index_offset_ack_0 : boolean;
  signal array_obj_ref_1098_index_offset_req_1 : boolean;
  signal array_obj_ref_1098_index_offset_ack_1 : boolean;
  signal array_obj_ref_1108_load_0_req_0 : boolean;
  signal array_obj_ref_1108_load_0_ack_0 : boolean;
  signal array_obj_ref_1108_load_0_req_1 : boolean;
  signal array_obj_ref_1108_load_0_ack_1 : boolean;
  signal array_obj_ref_1111_load_0_req_0 : boolean;
  signal array_obj_ref_1111_load_0_ack_0 : boolean;
  signal array_obj_ref_1111_load_0_req_1 : boolean;
  signal array_obj_ref_1111_load_0_ack_1 : boolean;
  signal type_cast_1113_inst_req_0 : boolean;
  signal type_cast_1113_inst_ack_0 : boolean;
  signal type_cast_1113_inst_req_1 : boolean;
  signal type_cast_1113_inst_ack_1 : boolean;
  signal array_obj_ref_1118_index_offset_req_0 : boolean;
  signal array_obj_ref_1118_index_offset_ack_0 : boolean;
  signal array_obj_ref_1118_index_offset_req_1 : boolean;
  signal array_obj_ref_1118_index_offset_ack_1 : boolean;
  signal array_obj_ref_1118_load_0_req_0 : boolean;
  signal array_obj_ref_1118_load_0_ack_0 : boolean;
  signal array_obj_ref_1118_load_0_req_1 : boolean;
  signal array_obj_ref_1118_load_0_ack_1 : boolean;
  signal array_obj_ref_1121_load_0_req_0 : boolean;
  signal array_obj_ref_1121_load_0_ack_0 : boolean;
  signal array_obj_ref_1121_load_0_req_1 : boolean;
  signal array_obj_ref_1121_load_0_ack_1 : boolean;
  signal type_cast_1123_inst_req_0 : boolean;
  signal type_cast_1123_inst_ack_0 : boolean;
  signal type_cast_1123_inst_req_1 : boolean;
  signal type_cast_1123_inst_ack_1 : boolean;
  signal array_obj_ref_1128_index_offset_req_0 : boolean;
  signal array_obj_ref_1128_index_offset_ack_0 : boolean;
  signal array_obj_ref_1128_index_offset_req_1 : boolean;
  signal array_obj_ref_1128_index_offset_ack_1 : boolean;
  signal array_obj_ref_1128_load_0_req_0 : boolean;
  signal array_obj_ref_1128_load_0_ack_0 : boolean;
  signal array_obj_ref_1128_load_0_req_1 : boolean;
  signal array_obj_ref_1128_load_0_ack_1 : boolean;
  signal array_obj_ref_1131_load_0_req_0 : boolean;
  signal array_obj_ref_1131_load_0_ack_0 : boolean;
  signal array_obj_ref_1131_load_0_req_1 : boolean;
  signal array_obj_ref_1131_load_0_ack_1 : boolean;
  signal type_cast_1133_inst_req_0 : boolean;
  signal type_cast_1133_inst_ack_0 : boolean;
  signal type_cast_1133_inst_req_1 : boolean;
  signal type_cast_1133_inst_ack_1 : boolean;
  signal array_obj_ref_1138_index_offset_req_0 : boolean;
  signal array_obj_ref_1138_index_offset_ack_0 : boolean;
  signal array_obj_ref_1138_index_offset_req_1 : boolean;
  signal array_obj_ref_1138_index_offset_ack_1 : boolean;
  signal array_obj_ref_1138_load_0_req_0 : boolean;
  signal array_obj_ref_1138_load_0_ack_0 : boolean;
  signal array_obj_ref_1138_load_0_req_1 : boolean;
  signal array_obj_ref_1138_load_0_ack_1 : boolean;
  signal array_obj_ref_1141_load_0_req_0 : boolean;
  signal array_obj_ref_1141_load_0_ack_0 : boolean;
  signal array_obj_ref_1141_load_0_req_1 : boolean;
  signal array_obj_ref_1141_load_0_ack_1 : boolean;
  signal type_cast_1143_inst_req_0 : boolean;
  signal type_cast_1143_inst_ack_0 : boolean;
  signal type_cast_1143_inst_req_1 : boolean;
  signal type_cast_1143_inst_ack_1 : boolean;
  signal type_cast_1149_inst_req_0 : boolean;
  signal type_cast_1149_inst_ack_0 : boolean;
  signal type_cast_1149_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_1 : boolean;
  signal type_cast_1155_inst_req_0 : boolean;
  signal type_cast_1155_inst_ack_0 : boolean;
  signal type_cast_1155_inst_req_1 : boolean;
  signal type_cast_1155_inst_ack_1 : boolean;
  signal type_cast_1161_inst_req_0 : boolean;
  signal type_cast_1161_inst_ack_0 : boolean;
  signal type_cast_1161_inst_req_1 : boolean;
  signal type_cast_1161_inst_ack_1 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal type_cast_1179_inst_req_0 : boolean;
  signal type_cast_1179_inst_ack_0 : boolean;
  signal type_cast_1179_inst_req_1 : boolean;
  signal type_cast_1179_inst_ack_1 : boolean;
  signal type_cast_1185_inst_req_0 : boolean;
  signal type_cast_1185_inst_ack_0 : boolean;
  signal type_cast_1185_inst_req_1 : boolean;
  signal type_cast_1185_inst_ack_1 : boolean;
  signal type_cast_1191_inst_req_0 : boolean;
  signal type_cast_1191_inst_ack_0 : boolean;
  signal type_cast_1191_inst_req_1 : boolean;
  signal type_cast_1191_inst_ack_1 : boolean;
  signal type_cast_1197_inst_req_0 : boolean;
  signal type_cast_1197_inst_ack_0 : boolean;
  signal type_cast_1197_inst_req_1 : boolean;
  signal type_cast_1197_inst_ack_1 : boolean;
  signal type_cast_1203_inst_req_0 : boolean;
  signal type_cast_1203_inst_ack_0 : boolean;
  signal type_cast_1203_inst_req_1 : boolean;
  signal type_cast_1203_inst_ack_1 : boolean;
  signal type_cast_1209_inst_req_0 : boolean;
  signal type_cast_1209_inst_ack_0 : boolean;
  signal type_cast_1209_inst_req_1 : boolean;
  signal type_cast_1209_inst_ack_1 : boolean;
  signal type_cast_1215_inst_req_0 : boolean;
  signal type_cast_1215_inst_ack_0 : boolean;
  signal type_cast_1215_inst_req_1 : boolean;
  signal type_cast_1215_inst_ack_1 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal type_cast_1227_inst_req_0 : boolean;
  signal type_cast_1227_inst_ack_0 : boolean;
  signal type_cast_1227_inst_req_1 : boolean;
  signal type_cast_1227_inst_ack_1 : boolean;
  signal type_cast_1233_inst_req_0 : boolean;
  signal type_cast_1233_inst_ack_0 : boolean;
  signal type_cast_1233_inst_req_1 : boolean;
  signal type_cast_1233_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "mainAcc2_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 13) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= I;
  I_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(10 downto 6) <= J;
  J_buffer <= in_buffer_data_out(10 downto 6);
  in_buffer_data_in(12 downto 11) <= col_to_be_replaced;
  col_to_be_replaced_buffer <= in_buffer_data_out(12 downto 11);
  in_buffer_data_in(tag_length + 12 downto 13) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 12 downto 13);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  mainAcc2_CP_4584_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "mainAcc2_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ofmap_pixel_buffer;
  ofmap_pixel <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mainAcc2_CP_4584_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= mainAcc2_CP_4584_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= mainAcc2_CP_4584_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,mainAcc2_CP_4584_start,"mainAcc2 cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,mainAcc2_CP_4584_symbol, "mainAcc2 cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  mainAcc2_CP_4584: Block -- control-path 
    signal mainAcc2_CP_4584_elements: BooleanArray(196 downto 0);
    -- 
  begin -- 
    mainAcc2_CP_4584_elements(0) <= mainAcc2_CP_4584_start;
    mainAcc2_CP_4584_symbol <= mainAcc2_CP_4584_elements(196);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	128 
    -- CP-element group 0: 	30 
    -- CP-element group 0: 	112 
    -- CP-element group 0: 	150 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	47 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	94 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	162 
    -- CP-element group 0: 	156 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	129 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	26 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	63 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	120 
    -- CP-element group 0: 	146 
    -- CP-element group 0: 	192 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	186 
    -- CP-element group 0: 	189 
    -- CP-element group 0: 	66 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	102 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	18 
    -- CP-element group 0: 	39 
    -- CP-element group 0: 	138 
    -- CP-element group 0: 	139 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	78 
    -- CP-element group 0: 	42 
    -- CP-element group 0: 	168 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	83 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	87 
    -- CP-element group 0: 	90 
    -- CP-element group 0: 	92 
    -- CP-element group 0: 	96 
    -- CP-element group 0: 	99 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	132 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	108 
    -- CP-element group 0: 	110 
    -- CP-element group 0: 	111 
    -- CP-element group 0: 	114 
    -- CP-element group 0: 	126 
    -- CP-element group 0: 	180 
    -- CP-element group 0: 	195 
    -- CP-element group 0: 	51 
    -- CP-element group 0: 	165 
    -- CP-element group 0: 	141 
    -- CP-element group 0: 	130 
    -- CP-element group 0: 	35 
    -- CP-element group 0: 	137 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	119 
    -- CP-element group 0: 	171 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	123 
    -- CP-element group 0: 	153 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	135 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	144 
    -- CP-element group 0: 	147 
    -- CP-element group 0: 	148 
    -- CP-element group 0: 	174 
    -- CP-element group 0: 	159 
    -- CP-element group 0: 	121 
    -- CP-element group 0: 	177 
    -- CP-element group 0: 	183 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	22 
    -- CP-element group 0: 	24 
    -- CP-element group 0:  members (485) 
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_resized_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_computed_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_computed_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_resized_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_resized_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_computed_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_resized_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_computed_1
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_start/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_complete/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_start/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_complete/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_start/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_complete/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_sample_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Update/cr
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_update_start_
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Update/$entry
      -- CP-element group 0: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Update/cr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1121_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1043_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1167_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1173_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1155_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1081_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1081_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1041_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1121_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1113_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_957_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_957_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_971_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_971_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1031_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1111_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1111_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1227_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1221_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1051_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1141_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1141_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_983_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_983_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_993_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1053_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1041_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1051_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_991_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_991_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1003_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1031_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1063_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1021_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1021_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1061_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1061_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1073_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1033_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1011_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1185_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1011_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1071_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1071_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1083_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1093_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1091_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1091_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1133_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1103_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1101_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1101_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1209_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1233_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1179_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1143_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1023_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1191_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1123_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1149_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_index_offset_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1131_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1131_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1197_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1161_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1203_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1215_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1001_load_0_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1001_load_0_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1013_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_6267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1121_load_0_req_1); -- 
    cr_5338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1043_inst_req_1); -- 
    cr_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1038_load_0_req_1); -- 
    req_4903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1008_index_offset_req_1); -- 
    cr_5053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1018_load_0_req_1); -- 
    req_5729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1078_index_offset_req_1); -- 
    req_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1028_index_offset_req_1); -- 
    cr_6574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1167_inst_req_1); -- 
    cr_6588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1173_inst_req_1); -- 
    req_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1018_index_offset_req_0); -- 
    cr_6546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1155_inst_req_1); -- 
    cr_5795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1081_load_0_req_1); -- 
    rr_5784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1081_load_0_req_0); -- 
    rr_5312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1041_load_0_req_0); -- 
    rr_6256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1121_load_0_req_0); -- 
    cr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1113_inst_req_1); -- 
    cr_6115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1108_load_0_req_1); -- 
    req_4597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_957_inst_req_0); -- 
    req_4602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_957_inst_req_1); -- 
    req_4611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_971_inst_req_0); -- 
    req_4616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_971_inst_req_1); -- 
    req_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1038_index_offset_req_1); -- 
    rr_5194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1031_load_0_req_0); -- 
    cr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1111_load_0_req_1); -- 
    rr_6138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1111_load_0_req_0); -- 
    cr_6714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1227_inst_req_1); -- 
    cr_6233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1118_load_0_req_1); -- 
    req_5375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1048_index_offset_req_1); -- 
    cr_6700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1221_inst_req_1); -- 
    cr_5407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1048_load_0_req_1); -- 
    rr_5430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1051_load_0_req_0); -- 
    cr_6503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1141_load_0_req_1); -- 
    rr_6492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1141_load_0_req_0); -- 
    req_4625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_983_inst_req_0); -- 
    req_4630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => MUX_983_inst_req_1); -- 
    cr_4748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_993_inst_req_1); -- 
    cr_4699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_988_load_0_req_1); -- 
    req_4898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1008_index_offset_req_0); -- 
    cr_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1053_inst_req_1); -- 
    cr_5323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1041_load_0_req_1); -- 
    cr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1051_load_0_req_1); -- 
    req_4662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_988_index_offset_req_0); -- 
    req_4667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_988_index_offset_req_1); -- 
    cr_4733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_991_load_0_req_1); -- 
    rr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_991_load_0_req_0); -- 
    cr_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1003_inst_req_1); -- 
    cr_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_998_load_0_req_1); -- 
    req_4780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_998_index_offset_req_0); -- 
    req_4785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_998_index_offset_req_1); -- 
    cr_5205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1031_load_0_req_1); -- 
    cr_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1063_inst_req_1); -- 
    cr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1058_load_0_req_1); -- 
    cr_5087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1021_load_0_req_1); -- 
    rr_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1021_load_0_req_0); -- 
    req_5493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1058_index_offset_req_1); -- 
    cr_5559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1061_load_0_req_1); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1061_load_0_req_0); -- 
    cr_5692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1073_inst_req_1); -- 
    cr_5643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1068_load_0_req_1); -- 
    cr_5220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1033_inst_req_1); -- 
    cr_5171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1028_load_0_req_1); -- 
    cr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1011_load_0_req_1); -- 
    req_5611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1068_index_offset_req_1); -- 
    cr_6616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1185_inst_req_1); -- 
    rr_4958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1011_load_0_req_0); -- 
    cr_5677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1071_load_0_req_1); -- 
    rr_5666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1071_load_0_req_0); -- 
    cr_5810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1083_inst_req_1); -- 
    cr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1078_load_0_req_1); -- 
    cr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1093_inst_req_1); -- 
    cr_5879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1088_load_0_req_1); -- 
    req_5847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1088_index_offset_req_1); -- 
    cr_5913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1091_load_0_req_1); -- 
    rr_5902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1091_load_0_req_0); -- 
    cr_6400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1133_inst_req_1); -- 
    cr_6046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1103_inst_req_1); -- 
    cr_5997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1098_load_0_req_1); -- 
    req_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1098_index_offset_req_1); -- 
    cr_6031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1101_load_0_req_1); -- 
    rr_6020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1101_load_0_req_0); -- 
    cr_6672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1209_inst_req_1); -- 
    cr_6728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1233_inst_req_1); -- 
    req_6083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1108_index_offset_req_1); -- 
    cr_6602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1179_inst_req_1); -- 
    cr_6518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1143_inst_req_1); -- 
    cr_6469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1138_load_0_req_1); -- 
    cr_6351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1128_load_0_req_1); -- 
    req_5021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1018_index_offset_req_1); -- 
    cr_5102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1023_inst_req_1); -- 
    cr_6630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1191_inst_req_1); -- 
    req_6437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1138_index_offset_req_1); -- 
    req_6201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1118_index_offset_req_1); -- 
    cr_6282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1123_inst_req_1); -- 
    cr_6532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1149_inst_req_1); -- 
    req_6319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1128_index_offset_req_1); -- 
    cr_6385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1131_load_0_req_1); -- 
    rr_6374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1131_load_0_req_0); -- 
    cr_6644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1197_inst_req_1); -- 
    cr_6560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1161_inst_req_1); -- 
    cr_6658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1203_inst_req_1); -- 
    cr_6686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1215_inst_req_1); -- 
    cr_4851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1001_load_0_req_1); -- 
    rr_4840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1001_load_0_req_0); -- 
    cr_4984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => type_cast_1013_inst_req_1); -- 
    cr_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(0), ack => array_obj_ref_1008_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_sample_completed_
      -- CP-element group 1: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_start/$exit
      -- CP-element group 1: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_start/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_957_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_957_inst_ack_0, ack => mainAcc2_CP_4584_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	44 
    -- CP-element group 2: 	53 
    -- CP-element group 2: 	62 
    -- CP-element group 2: 	71 
    -- CP-element group 2:  members (55) 
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_update_completed_
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_complete/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/MUX_957_complete/ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_resized_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_computed_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_resized_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_computed_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_resized_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_computed_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Sample/req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_resized_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_scaled_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_computed_1
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_resize_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_resize_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_resize_1/index_resize_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_resize_1/index_resize_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_scale_1/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_scale_1/$exit
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_scale_1/scale_rename_req
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_index_scale_1/scale_rename_ack
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_957_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_957_inst_ack_1, ack => mainAcc2_CP_4584_elements(2)); -- 
    req_5370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(2), ack => array_obj_ref_1048_index_offset_req_0); -- 
    req_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(2), ack => array_obj_ref_1058_index_offset_req_0); -- 
    req_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(2), ack => array_obj_ref_1028_index_offset_req_0); -- 
    req_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(2), ack => array_obj_ref_1038_index_offset_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_sample_completed_
      -- CP-element group 3: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_start/$exit
      -- CP-element group 3: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_start/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_971_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_971_inst_ack_0, ack => mainAcc2_CP_4584_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	89 
    -- CP-element group 4: 	80 
    -- CP-element group 4: 	98 
    -- CP-element group 4: 	107 
    -- CP-element group 4:  members (55) 
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_update_completed_
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_complete/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/MUX_971_complete/ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_resized_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_computed_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_resized_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_computed_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_resized_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_computed_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Sample/req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_resized_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_scaled_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_computed_1
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_resize_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_resize_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_resize_1/index_resize_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_resize_1/index_resize_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_scale_1/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_scale_1/$exit
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_scale_1/scale_rename_req
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_index_scale_1/scale_rename_ack
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_971_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_971_inst_ack_1, ack => mainAcc2_CP_4584_elements(4)); -- 
    req_5606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(4), ack => array_obj_ref_1068_index_offset_req_0); -- 
    req_5724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(4), ack => array_obj_ref_1078_index_offset_req_0); -- 
    req_5960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(4), ack => array_obj_ref_1098_index_offset_req_0); -- 
    req_5842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(4), ack => array_obj_ref_1088_index_offset_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_sample_completed_
      -- CP-element group 5: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_start/$exit
      -- CP-element group 5: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_start/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_983_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_983_inst_ack_0, ack => mainAcc2_CP_4584_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	143 
    -- CP-element group 6: 	125 
    -- CP-element group 6: 	134 
    -- CP-element group 6: 	116 
    -- CP-element group 6:  members (55) 
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_update_completed_
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_complete/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/MUX_983_complete/ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_computed_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_index_resized_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_resized_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_computed_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_resized_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_computed_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Sample/req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_resized_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_scaled_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_computed_1
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_resize_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_resize_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_resize_1/index_resize_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_resize_1/index_resize_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_scale_1/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_scale_1/$exit
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_scale_1/scale_rename_req
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_index_scale_1/scale_rename_ack
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Sample/$entry
      -- CP-element group 6: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Sample/req
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:MUX_983_inst_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_index_offset_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_index_offset_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_983_inst_ack_1, ack => mainAcc2_CP_4584_elements(6)); -- 
    req_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(6), ack => array_obj_ref_1118_index_offset_req_0); -- 
    req_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(6), ack => array_obj_ref_1108_index_offset_req_0); -- 
    req_6432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(6), ack => array_obj_ref_1138_index_offset_req_0); -- 
    req_6314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(6), ack => array_obj_ref_1128_index_offset_req_0); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	11 
    -- CP-element group 7: 	13 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	14 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Sample/$entry
      -- CP-element group 7: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Sample/rr
      -- CP-element group 7: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_sample_start_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_993_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(7), ack => type_cast_993_inst_req_0); -- 
    mainAcc2_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "mainAcc2_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(11) & mainAcc2_CP_4584_elements(13);
      gj_mainAcc2_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	196 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Sample/ack
      -- CP-element group 8: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_sample_complete
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_988_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (18) 
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_word_addrgen/$exit
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_sample_start_
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_word_addrgen/root_register_ack
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_word_addrgen/root_register_req
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/$entry
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_word_address_calculated
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Update/$exit
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_final_index_sum_regn_Update/ack
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_base_plus_offset/$entry
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/word_0/$entry
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_base_plus_offset/$exit
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/word_0/rr
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_base_plus_offset/sum_rename_req
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_base_plus_offset/sum_rename_ack
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_root_address_calculated
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_offset_calculated
      -- CP-element group 9: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_word_addrgen/$entry
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_988_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(9)); -- 
    rr_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(9), ack => array_obj_ref_988_load_0_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_sample_completed_
      -- CP-element group 10: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/$exit
      -- CP-element group 10: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/$exit
      -- CP-element group 10: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_988_load_0_ack_0, ack => mainAcc2_CP_4584_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	7 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/array_obj_ref_988_Merge/$exit
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_update_completed_
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/array_obj_ref_988_Merge/merge_ack
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/array_obj_ref_988_Merge/merge_req
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/word_0/ca
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/array_obj_ref_988_Merge/$entry
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/word_access_complete/$exit
      -- CP-element group 11: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_988_Update/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_988_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_988_load_0_ack_1, ack => mainAcc2_CP_4584_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_sample_completed_
      -- CP-element group 12: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/$exit
      -- CP-element group 12: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/word_0/$exit
      -- CP-element group 12: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_991_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_991_load_0_ack_0, ack => mainAcc2_CP_4584_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	7 
    -- CP-element group 13:  members (9) 
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/word_0/$exit
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_update_completed_
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/array_obj_ref_991_Merge/$entry
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/$exit
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/array_obj_ref_991_Merge/merge_ack
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/word_0/ca
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/array_obj_ref_991_Merge/$exit
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/array_obj_ref_991_Merge/merge_req
      -- CP-element group 13: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_991_Update/word_access_complete/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_991_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_991_load_0_ack_1, ack => mainAcc2_CP_4584_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	7 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Sample/$exit
      -- CP-element group 14: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Sample/ra
      -- CP-element group 14: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_sample_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_993_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_993_inst_ack_0, ack => mainAcc2_CP_4584_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	154 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Update/$exit
      -- CP-element group 15: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_Update/ca
      -- CP-element group 15: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_993_update_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_993_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_993_inst_ack_1, ack => mainAcc2_CP_4584_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	22 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Sample/rr
      -- CP-element group 16: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_sample_start_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1003_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(16), ack => type_cast_1003_inst_req_0); -- 
    mainAcc2_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(20) & mainAcc2_CP_4584_elements(22);
      gj_mainAcc2_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	196 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Sample/ack
      -- CP-element group 17: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Sample/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	0 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (18) 
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_offset_calculated
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_word_address_calculated
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/$entry
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/word_0/rr
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_root_address_calculated
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_word_addrgen/$entry
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/word_0/$entry
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_word_addrgen/$exit
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/$entry
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_sample_start_
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_word_addrgen/root_register_req
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_word_addrgen/root_register_ack
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_base_plus_offset/$exit
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_base_plus_offset/$entry
      -- CP-element group 18: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_final_index_sum_regn_Update/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(18)); -- 
    rr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(18), ack => array_obj_ref_998_load_0_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_sample_completed_
      -- CP-element group 19: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Sample/word_access_start/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_load_0_ack_0, ack => mainAcc2_CP_4584_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/$exit
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_update_completed_
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/word_access_complete/$exit
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/array_obj_ref_998_Merge/$entry
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/array_obj_ref_998_Merge/$exit
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/array_obj_ref_998_Merge/merge_req
      -- CP-element group 20: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_998_Update/array_obj_ref_998_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_998_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_load_0_ack_1, ack => mainAcc2_CP_4584_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/$exit
      -- CP-element group 21: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/$exit
      -- CP-element group 21: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Sample/word_access_start/word_0/ra
      -- CP-element group 21: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_sample_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1001_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1001_load_0_ack_0, ack => mainAcc2_CP_4584_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	0 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	16 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/array_obj_ref_1001_Merge/merge_ack
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/array_obj_ref_1001_Merge/merge_req
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/$exit
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/$exit
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/array_obj_ref_1001_Merge/$exit
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_update_completed_
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/array_obj_ref_1001_Merge/$entry
      -- CP-element group 22: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1001_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1001_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1001_load_0_ack_1, ack => mainAcc2_CP_4584_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Sample/$exit
      -- CP-element group 23: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_sample_completed_
      -- CP-element group 23: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1003_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1003_inst_ack_0, ack => mainAcc2_CP_4584_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	160 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Update/ca
      -- CP-element group 24: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_update_completed_
      -- CP-element group 24: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1003_Update/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1003_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1003_inst_ack_1, ack => mainAcc2_CP_4584_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	31 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	32 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_sample_start_
      -- CP-element group 25: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Sample/$entry
      -- CP-element group 25: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1013_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(25), ack => type_cast_1013_inst_req_0); -- 
    mainAcc2_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(31) & mainAcc2_CP_4584_elements(29);
      gj_mainAcc2_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	0 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	196 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_sample_complete
      -- CP-element group 26: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Sample/ack
      -- CP-element group 26: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Sample/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (18) 
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_word_addrgen/$entry
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_base_plus_offset/$entry
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_word_addrgen/root_register_ack
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_root_address_calculated
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/word_0/rr
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/$entry
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Update/ack
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_offset_calculated
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_base_plus_offset/$exit
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_base_plus_offset/sum_rename_req
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_word_addrgen/$exit
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_word_addrgen/root_register_req
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/word_0/$entry
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_word_address_calculated
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_base_plus_offset/sum_rename_ack
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_sample_start_
      -- CP-element group 27: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_final_index_sum_regn_Update/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_4904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(27)); -- 
    rr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(27), ack => array_obj_ref_1008_load_0_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (5) 
      -- CP-element group 28: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_sample_completed_
      -- CP-element group 28: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/word_0/ra
      -- CP-element group 28: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/$exit
      -- CP-element group 28: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/$exit
      -- CP-element group 28: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Sample/word_access_start/word_0/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_load_0_ack_0, ack => mainAcc2_CP_4584_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/array_obj_ref_1008_Merge/$exit
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/$exit
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_update_completed_
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/word_0/$exit
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/word_access_complete/word_0/ca
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/$exit
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/array_obj_ref_1008_Merge/$entry
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/array_obj_ref_1008_Merge/merge_req
      -- CP-element group 29: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1008_Update/array_obj_ref_1008_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1008_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1008_load_0_ack_1, ack => mainAcc2_CP_4584_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	0 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/$exit
      -- CP-element group 30: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_sample_completed_
      -- CP-element group 30: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/word_0/$exit
      -- CP-element group 30: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/$exit
      -- CP-element group 30: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1011_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1011_load_0_ack_0, ack => mainAcc2_CP_4584_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	25 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_update_completed_
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/$exit
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/array_obj_ref_1011_Merge/$entry
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/array_obj_ref_1011_Merge/$exit
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/array_obj_ref_1011_Merge/merge_req
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/array_obj_ref_1011_Merge/merge_ack
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/word_0/ca
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/$exit
      -- CP-element group 31: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1011_Update/word_access_complete/word_0/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1011_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1011_load_0_ack_1, ack => mainAcc2_CP_4584_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	25 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_sample_completed_
      -- CP-element group 32: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Sample/ra
      -- CP-element group 32: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Sample/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1013_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_0, ack => mainAcc2_CP_4584_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	166 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_update_completed_
      -- CP-element group 33: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Update/ca
      -- CP-element group 33: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1013_Update/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1013_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_4985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_1, ack => mainAcc2_CP_4584_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	38 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	41 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_sample_start_
      -- CP-element group 34: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1023_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(34), ack => type_cast_1023_inst_req_0); -- 
    mainAcc2_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(40) & mainAcc2_CP_4584_elements(38);
      gj_mainAcc2_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	196 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_sample_complete
      -- CP-element group 35: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1018_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(35)); -- 
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (18) 
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_root_address_calculated
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_offset_calculated
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_sample_start_
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_word_address_calculated
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Update/$exit
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_final_index_sum_regn_Update/ack
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_base_plus_offset/$entry
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_base_plus_offset/$exit
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_base_plus_offset/sum_rename_req
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_base_plus_offset/sum_rename_ack
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_word_addrgen/$entry
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_word_addrgen/$exit
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_word_addrgen/root_register_req
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_word_addrgen/root_register_ack
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/$entry
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1018_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(36)); -- 
    rr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(36), ack => array_obj_ref_1018_load_0_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_sample_completed_
      -- CP-element group 37: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/$exit
      -- CP-element group 37: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/$exit
      -- CP-element group 37: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/word_0/$exit
      -- CP-element group 37: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1018_load_0_ack_0, ack => mainAcc2_CP_4584_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	34 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_update_completed_
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/$exit
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/$exit
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/word_access_complete/word_0/ca
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/array_obj_ref_1018_Merge/$entry
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/array_obj_ref_1018_Merge/$exit
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/array_obj_ref_1018_Merge/merge_req
      -- CP-element group 38: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1018_Update/array_obj_ref_1018_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1018_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1018_load_0_ack_1, ack => mainAcc2_CP_4584_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	0 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_sample_completed_
      -- CP-element group 39: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/$exit
      -- CP-element group 39: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/$exit
      -- CP-element group 39: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1021_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_load_0_ack_0, ack => mainAcc2_CP_4584_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	34 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_update_completed_
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/$exit
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/$exit
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/word_0/$exit
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/word_access_complete/word_0/ca
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/array_obj_ref_1021_Merge/$entry
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/array_obj_ref_1021_Merge/$exit
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/array_obj_ref_1021_Merge/merge_req
      -- CP-element group 40: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1021_Update/array_obj_ref_1021_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1021_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_load_0_ack_1, ack => mainAcc2_CP_4584_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_sample_completed_
      -- CP-element group 41: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Sample/$exit
      -- CP-element group 41: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1023_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1023_inst_ack_0, ack => mainAcc2_CP_4584_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	0 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	172 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_update_completed_
      -- CP-element group 42: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Update/$exit
      -- CP-element group 42: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1023_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1023_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1023_inst_ack_1, ack => mainAcc2_CP_4584_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	49 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	50 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_sample_start_
      -- CP-element group 43: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Sample/$entry
      -- CP-element group 43: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1033_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(43), ack => type_cast_1033_inst_req_0); -- 
    mainAcc2_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(47) & mainAcc2_CP_4584_elements(49);
      gj_mainAcc2_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	2 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	196 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_sample_complete
      -- CP-element group 44: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Sample/$exit
      -- CP-element group 44: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (18) 
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_sample_start_
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_word_address_calculated
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_root_address_calculated
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_offset_calculated
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Update/$exit
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_final_index_sum_regn_Update/ack
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_base_plus_offset/$entry
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_base_plus_offset/$exit
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_word_addrgen/$entry
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_word_addrgen/$exit
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_word_addrgen/root_register_req
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_word_addrgen/root_register_ack
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/$entry
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/$entry
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(45)); -- 
    rr_5160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(45), ack => array_obj_ref_1028_load_0_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_sample_completed_
      -- CP-element group 46: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_load_0_ack_0, ack => mainAcc2_CP_4584_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	0 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	43 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_update_completed_
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/$exit
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/array_obj_ref_1028_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/array_obj_ref_1028_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/array_obj_ref_1028_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1028_Update/array_obj_ref_1028_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1028_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_load_0_ack_1, ack => mainAcc2_CP_4584_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_sample_completed_
      -- CP-element group 48: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/$exit
      -- CP-element group 48: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/$exit
      -- CP-element group 48: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/word_0/$exit
      -- CP-element group 48: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1031_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1031_load_0_ack_0, ack => mainAcc2_CP_4584_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	43 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_update_completed_
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/$exit
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/$exit
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/word_0/$exit
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/word_access_complete/word_0/ca
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/array_obj_ref_1031_Merge/$entry
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/array_obj_ref_1031_Merge/$exit
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/array_obj_ref_1031_Merge/merge_req
      -- CP-element group 49: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1031_Update/array_obj_ref_1031_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1031_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1031_load_0_ack_1, ack => mainAcc2_CP_4584_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	43 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_sample_completed_
      -- CP-element group 50: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1033_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_0, ack => mainAcc2_CP_4584_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	0 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	154 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_update_completed_
      -- CP-element group 51: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Update/$exit
      -- CP-element group 51: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1033_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1033_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_1, ack => mainAcc2_CP_4584_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	58 
    -- CP-element group 52: 	56 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	59 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_sample_start_
      -- CP-element group 52: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1043_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(52), ack => type_cast_1043_inst_req_0); -- 
    mainAcc2_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(58) & mainAcc2_CP_4584_elements(56);
      gj_mainAcc2_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	2 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	196 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_sample_complete
      -- CP-element group 53: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Sample/$exit
      -- CP-element group 53: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (18) 
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_sample_start_
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_word_address_calculated
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_root_address_calculated
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_offset_calculated
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Update/$exit
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_final_index_sum_regn_Update/ack
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_base_plus_offset/$entry
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_base_plus_offset/$exit
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_word_addrgen/$entry
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_word_addrgen/$exit
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_word_addrgen/root_register_req
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_word_addrgen/root_register_ack
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/$entry
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/$entry
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/word_0/$entry
      -- CP-element group 54: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(54)); -- 
    rr_5278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(54), ack => array_obj_ref_1038_load_0_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_sample_completed_
      -- CP-element group 55: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/$exit
      -- CP-element group 55: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/$exit
      -- CP-element group 55: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/word_0/$exit
      -- CP-element group 55: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_load_0_ack_0, ack => mainAcc2_CP_4584_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	52 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_update_completed_
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/$exit
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/$exit
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/word_0/$exit
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/word_access_complete/word_0/ca
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/array_obj_ref_1038_Merge/$entry
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/array_obj_ref_1038_Merge/$exit
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/array_obj_ref_1038_Merge/merge_req
      -- CP-element group 56: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1038_Update/array_obj_ref_1038_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1038_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1038_load_0_ack_1, ack => mainAcc2_CP_4584_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_sample_completed_
      -- CP-element group 57: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/$exit
      -- CP-element group 57: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/$exit
      -- CP-element group 57: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/word_0/$exit
      -- CP-element group 57: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1041_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1041_load_0_ack_0, ack => mainAcc2_CP_4584_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	52 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_update_completed_
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/$exit
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/$exit
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/word_0/$exit
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/word_access_complete/word_0/ca
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/array_obj_ref_1041_Merge/$entry
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/array_obj_ref_1041_Merge/$exit
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/array_obj_ref_1041_Merge/merge_req
      -- CP-element group 58: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1041_Update/array_obj_ref_1041_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1041_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1041_load_0_ack_1, ack => mainAcc2_CP_4584_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	52 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_sample_completed_
      -- CP-element group 59: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Sample/$exit
      -- CP-element group 59: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1043_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1043_inst_ack_0, ack => mainAcc2_CP_4584_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	160 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_update_completed_
      -- CP-element group 60: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Update/$exit
      -- CP-element group 60: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1043_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1043_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1043_inst_ack_1, ack => mainAcc2_CP_4584_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	67 
    -- CP-element group 61: 	65 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	68 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_sample_start_
      -- CP-element group 61: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Sample/$entry
      -- CP-element group 61: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1053_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(61), ack => type_cast_1053_inst_req_0); -- 
    mainAcc2_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(67) & mainAcc2_CP_4584_elements(65);
      gj_mainAcc2_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	2 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	196 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_sample_complete
      -- CP-element group 62: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	0 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_sample_start_
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_word_address_calculated
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_root_address_calculated
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_offset_calculated
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Update/$exit
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_final_index_sum_regn_Update/ack
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_base_plus_offset/$entry
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_base_plus_offset/$exit
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_word_addrgen/$entry
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_word_addrgen/$exit
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_word_addrgen/root_register_req
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_word_addrgen/root_register_ack
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/$entry
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/$entry
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(63)); -- 
    rr_5396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(63), ack => array_obj_ref_1048_load_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_sample_completed_
      -- CP-element group 64: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/$exit
      -- CP-element group 64: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_load_0_ack_0, ack => mainAcc2_CP_4584_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	61 
    -- CP-element group 65:  members (9) 
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_update_completed_
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/$exit
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/$exit
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/array_obj_ref_1048_Merge/$entry
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/array_obj_ref_1048_Merge/$exit
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/array_obj_ref_1048_Merge/merge_req
      -- CP-element group 65: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1048_Update/array_obj_ref_1048_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1048_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_load_0_ack_1, ack => mainAcc2_CP_4584_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	0 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_sample_completed_
      -- CP-element group 66: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/$exit
      -- CP-element group 66: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/word_0/$exit
      -- CP-element group 66: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1051_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1051_load_0_ack_0, ack => mainAcc2_CP_4584_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	61 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_update_completed_
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/$exit
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/$exit
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/word_0/$exit
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/word_access_complete/word_0/ca
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/array_obj_ref_1051_Merge/$entry
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/array_obj_ref_1051_Merge/$exit
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/array_obj_ref_1051_Merge/merge_req
      -- CP-element group 67: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1051_Update/array_obj_ref_1051_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1051_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1051_load_0_ack_1, ack => mainAcc2_CP_4584_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	61 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_sample_completed_
      -- CP-element group 68: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Sample/$exit
      -- CP-element group 68: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1053_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1053_inst_ack_0, ack => mainAcc2_CP_4584_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	166 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_update_completed_
      -- CP-element group 69: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Update/$exit
      -- CP-element group 69: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1053_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1053_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1053_inst_ack_1, ack => mainAcc2_CP_4584_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	74 
    -- CP-element group 70: 	76 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	77 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_sample_start_
      -- CP-element group 70: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Sample/$entry
      -- CP-element group 70: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(70) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1063_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(70), ack => type_cast_1063_inst_req_0); -- 
    mainAcc2_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(74) & mainAcc2_CP_4584_elements(76);
      gj_mainAcc2_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	2 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	196 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_sample_complete
      -- CP-element group 71: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Sample/$exit
      -- CP-element group 71: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (18) 
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_sample_start_
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_word_address_calculated
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_root_address_calculated
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_offset_calculated
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Update/$exit
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_final_index_sum_regn_Update/ack
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_base_plus_offset/$entry
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_base_plus_offset/$exit
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_word_addrgen/$entry
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_word_addrgen/$exit
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_word_addrgen/root_register_req
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_word_addrgen/root_register_ack
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/$entry
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(72)); -- 
    rr_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(72), ack => array_obj_ref_1058_load_0_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_sample_completed_
      -- CP-element group 73: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/$exit
      -- CP-element group 73: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/$exit
      -- CP-element group 73: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/word_0/$exit
      -- CP-element group 73: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_load_0_ack_0, ack => mainAcc2_CP_4584_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	70 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_update_completed_
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/$exit
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/$exit
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/word_0/$exit
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/word_access_complete/word_0/ca
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/array_obj_ref_1058_Merge/$entry
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/array_obj_ref_1058_Merge/$exit
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/array_obj_ref_1058_Merge/merge_req
      -- CP-element group 74: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1058_Update/array_obj_ref_1058_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1058_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_load_0_ack_1, ack => mainAcc2_CP_4584_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_sample_completed_
      -- CP-element group 75: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/$exit
      -- CP-element group 75: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/$exit
      -- CP-element group 75: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/word_0/$exit
      -- CP-element group 75: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1061_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1061_load_0_ack_0, ack => mainAcc2_CP_4584_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	70 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_update_completed_
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/$exit
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/$exit
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/word_0/$exit
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/word_access_complete/word_0/ca
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/array_obj_ref_1061_Merge/$entry
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/array_obj_ref_1061_Merge/$exit
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/array_obj_ref_1061_Merge/merge_req
      -- CP-element group 76: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1061_Update/array_obj_ref_1061_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1061_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1061_load_0_ack_1, ack => mainAcc2_CP_4584_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	70 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_sample_completed_
      -- CP-element group 77: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Sample/$exit
      -- CP-element group 77: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1063_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1063_inst_ack_0, ack => mainAcc2_CP_4584_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	0 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	172 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_update_completed_
      -- CP-element group 78: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Update/$exit
      -- CP-element group 78: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1063_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(78) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1063_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1063_inst_ack_1, ack => mainAcc2_CP_4584_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	85 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_sample_start_
      -- CP-element group 79: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Sample/$entry
      -- CP-element group 79: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1073_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(79), ack => type_cast_1073_inst_req_0); -- 
    mainAcc2_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(83) & mainAcc2_CP_4584_elements(85);
      gj_mainAcc2_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	4 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	196 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_sample_complete
      -- CP-element group 80: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Sample/$exit
      -- CP-element group 80: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1068_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (18) 
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_sample_start_
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_word_address_calculated
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_root_address_calculated
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_offset_calculated
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Update/$exit
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_final_index_sum_regn_Update/ack
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_base_plus_offset/$entry
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_base_plus_offset/$exit
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_base_plus_offset/sum_rename_req
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_base_plus_offset/sum_rename_ack
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_word_addrgen/$entry
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_word_addrgen/$exit
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_word_addrgen/root_register_req
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_word_addrgen/root_register_ack
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/$entry
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/$entry
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/word_0/$entry
      -- CP-element group 81: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(81) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1068_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(81)); -- 
    rr_5632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(81), ack => array_obj_ref_1068_load_0_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_sample_completed_
      -- CP-element group 82: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/$exit
      -- CP-element group 82: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(82) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1068_load_0_ack_0, ack => mainAcc2_CP_4584_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_update_completed_
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/$exit
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/$exit
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/array_obj_ref_1068_Merge/$entry
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/array_obj_ref_1068_Merge/$exit
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/array_obj_ref_1068_Merge/merge_req
      -- CP-element group 83: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1068_Update/array_obj_ref_1068_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(83) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1068_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1068_load_0_ack_1, ack => mainAcc2_CP_4584_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_sample_completed_
      -- CP-element group 84: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/$exit
      -- CP-element group 84: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/$exit
      -- CP-element group 84: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(84) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1071_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1071_load_0_ack_0, ack => mainAcc2_CP_4584_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	79 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_update_completed_
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/$exit
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/$exit
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/array_obj_ref_1071_Merge/$entry
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/array_obj_ref_1071_Merge/$exit
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/array_obj_ref_1071_Merge/merge_req
      -- CP-element group 85: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1071_Update/array_obj_ref_1071_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1071_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1071_load_0_ack_1, ack => mainAcc2_CP_4584_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	79 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_sample_completed_
      -- CP-element group 86: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1073_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_0, ack => mainAcc2_CP_4584_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	0 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	151 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_update_completed_
      -- CP-element group 87: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Update/$exit
      -- CP-element group 87: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1073_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1073_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_1, ack => mainAcc2_CP_4584_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	94 
    -- CP-element group 88: 	92 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	95 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_sample_start_
      -- CP-element group 88: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1083_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(88), ack => type_cast_1083_inst_req_0); -- 
    mainAcc2_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(94) & mainAcc2_CP_4584_elements(92);
      gj_mainAcc2_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	4 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	196 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_sample_complete
      -- CP-element group 89: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Sample/$exit
      -- CP-element group 89: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	0 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (18) 
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_sample_start_
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_word_address_calculated
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_root_address_calculated
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_offset_calculated
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Update/$exit
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_final_index_sum_regn_Update/ack
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_base_plus_offset/$entry
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_base_plus_offset/$exit
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_word_addrgen/$entry
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_word_addrgen/$exit
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_word_addrgen/root_register_req
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_word_addrgen/root_register_ack
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/$entry
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/$entry
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/word_0/$entry
      -- CP-element group 90: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(90)); -- 
    rr_5750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(90), ack => array_obj_ref_1078_load_0_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_sample_completed_
      -- CP-element group 91: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/$exit
      -- CP-element group 91: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_load_0_ack_0, ack => mainAcc2_CP_4584_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	0 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	88 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_update_completed_
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/$exit
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/$exit
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/word_access_complete/word_0/ca
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/array_obj_ref_1078_Merge/$entry
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/array_obj_ref_1078_Merge/$exit
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/array_obj_ref_1078_Merge/merge_req
      -- CP-element group 92: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1078_Update/array_obj_ref_1078_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1078_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_load_0_ack_1, ack => mainAcc2_CP_4584_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_sample_completed_
      -- CP-element group 93: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/$exit
      -- CP-element group 93: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1081_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1081_load_0_ack_0, ack => mainAcc2_CP_4584_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	0 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	88 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_update_completed_
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/$exit
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/$exit
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/array_obj_ref_1081_Merge/$entry
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/array_obj_ref_1081_Merge/$exit
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/array_obj_ref_1081_Merge/merge_req
      -- CP-element group 94: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1081_Update/array_obj_ref_1081_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1081_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1081_load_0_ack_1, ack => mainAcc2_CP_4584_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	88 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_sample_completed_
      -- CP-element group 95: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Sample/$exit
      -- CP-element group 95: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1083_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_0, ack => mainAcc2_CP_4584_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	0 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	157 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_update_completed_
      -- CP-element group 96: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Update/$exit
      -- CP-element group 96: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1083_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1083_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_1, ack => mainAcc2_CP_4584_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	103 
    -- CP-element group 97: 	101 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_sample_start_
      -- CP-element group 97: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Sample/$entry
      -- CP-element group 97: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1093_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(97), ack => type_cast_1093_inst_req_0); -- 
    mainAcc2_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "mainAcc2_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(103) & mainAcc2_CP_4584_elements(101);
      gj_mainAcc2_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	4 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	196 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_sample_complete
      -- CP-element group 98: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	0 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (18) 
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_sample_start_
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_word_address_calculated
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_root_address_calculated
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_offset_calculated
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Update/$exit
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_final_index_sum_regn_Update/ack
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_base_plus_offset/$entry
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_base_plus_offset/$exit
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_base_plus_offset/sum_rename_req
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_base_plus_offset/sum_rename_ack
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_word_addrgen/$entry
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_word_addrgen/$exit
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_word_addrgen/root_register_req
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_word_addrgen/root_register_ack
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/$entry
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/$entry
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/word_0/$entry
      -- CP-element group 99: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(99)); -- 
    rr_5868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(99), ack => array_obj_ref_1088_load_0_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_sample_completed_
      -- CP-element group 100: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/$exit
      -- CP-element group 100: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/$exit
      -- CP-element group 100: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/word_0/$exit
      -- CP-element group 100: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_load_0_ack_0, ack => mainAcc2_CP_4584_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	97 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_update_completed_
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/$exit
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/$exit
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/word_0/$exit
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/word_access_complete/word_0/ca
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/array_obj_ref_1088_Merge/$entry
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/array_obj_ref_1088_Merge/$exit
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/array_obj_ref_1088_Merge/merge_req
      -- CP-element group 101: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1088_Update/array_obj_ref_1088_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1088_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_load_0_ack_1, ack => mainAcc2_CP_4584_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	0 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_sample_completed_
      -- CP-element group 102: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/$exit
      -- CP-element group 102: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1091_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_load_0_ack_0, ack => mainAcc2_CP_4584_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	97 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_update_completed_
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/$exit
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/$exit
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/$entry
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/$exit
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/merge_req
      -- CP-element group 103: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1091_Update/array_obj_ref_1091_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1091_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_load_0_ack_1, ack => mainAcc2_CP_4584_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	97 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_sample_completed_
      -- CP-element group 104: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Sample/$exit
      -- CP-element group 104: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1093_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1093_inst_ack_0, ack => mainAcc2_CP_4584_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	163 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_update_completed_
      -- CP-element group 105: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Update/$exit
      -- CP-element group 105: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1093_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1093_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1093_inst_ack_1, ack => mainAcc2_CP_4584_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	112 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	113 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Sample/rr
      -- CP-element group 106: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Sample/$entry
      -- CP-element group 106: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_sample_start_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1103_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(106), ack => type_cast_1103_inst_req_0); -- 
    mainAcc2_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(112) & mainAcc2_CP_4584_elements(110);
      gj_mainAcc2_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	4 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	196 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_sample_complete
      -- CP-element group 107: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Sample/$exit
      -- CP-element group 107: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	0 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (18) 
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/word_0/rr
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_word_addrgen/root_register_ack
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/$entry
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_word_addrgen/root_register_req
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_word_addrgen/$exit
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_word_addrgen/$entry
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_sample_start_
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_word_address_calculated
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_root_address_calculated
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_offset_calculated
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Update/$exit
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_final_index_sum_regn_Update/ack
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_base_plus_offset/$entry
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_base_plus_offset/$exit
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_base_plus_offset/sum_rename_req
      -- CP-element group 108: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_base_plus_offset/sum_rename_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(108)); -- 
    rr_5986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(108), ack => array_obj_ref_1098_load_0_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/$exit
      -- CP-element group 109: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/$exit
      -- CP-element group 109: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_sample_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_5987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_load_0_ack_0, ack => mainAcc2_CP_4584_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	0 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/$exit
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/$exit
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/array_obj_ref_1098_Merge/merge_ack
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/array_obj_ref_1098_Merge/merge_req
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/array_obj_ref_1098_Merge/$exit
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/array_obj_ref_1098_Merge/$entry
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1098_update_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1098_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_5998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_load_0_ack_1, ack => mainAcc2_CP_4584_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	0 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/word_0/ra
      -- CP-element group 111: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/word_access_start/$exit
      -- CP-element group 111: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Sample/$exit
      -- CP-element group 111: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_sample_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1101_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1101_load_0_ack_0, ack => mainAcc2_CP_4584_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	0 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	106 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/array_obj_ref_1101_Merge/merge_ack
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/array_obj_ref_1101_Merge/merge_req
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/array_obj_ref_1101_Merge/$exit
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/array_obj_ref_1101_Merge/$entry
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/word_access_complete/$exit
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_Update/$exit
      -- CP-element group 112: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1101_update_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1101_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1101_load_0_ack_1, ack => mainAcc2_CP_4584_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	106 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Sample/ra
      -- CP-element group 113: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Sample/$exit
      -- CP-element group 113: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_sample_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1103_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1103_inst_ack_0, ack => mainAcc2_CP_4584_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	0 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	169 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Update/$exit
      -- CP-element group 114: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_Update/ca
      -- CP-element group 114: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1103_update_completed_
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1103_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1103_inst_ack_1, ack => mainAcc2_CP_4584_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	119 
    -- CP-element group 115: 	121 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_sample_start_
      -- CP-element group 115: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Sample/$entry
      -- CP-element group 115: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1113_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(115), ack => type_cast_1113_inst_req_0); -- 
    mainAcc2_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(119) & mainAcc2_CP_4584_elements(121);
      gj_mainAcc2_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	6 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	196 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_sample_complete
      -- CP-element group 116: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Sample/$exit
      -- CP-element group 116: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1108_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (18) 
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_sample_start_
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Update/$exit
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_final_index_sum_regn_Update/ack
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_offset_calculated
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_root_address_calculated
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_word_address_calculated
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_base_plus_offset/$entry
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_base_plus_offset/$exit
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_base_plus_offset/sum_rename_req
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_base_plus_offset/sum_rename_ack
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_word_addrgen/$entry
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_word_addrgen/$exit
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_word_addrgen/root_register_req
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_word_addrgen/root_register_ack
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/$entry
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/$entry
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1108_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(117)); -- 
    rr_6104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(117), ack => array_obj_ref_1108_load_0_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_sample_completed_
      -- CP-element group 118: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/$exit
      -- CP-element group 118: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/word_0/$exit
      -- CP-element group 118: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1108_load_0_ack_0, ack => mainAcc2_CP_4584_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	0 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	115 
    -- CP-element group 119:  members (9) 
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_update_completed_
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/$exit
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/$exit
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/word_0/$exit
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/word_access_complete/word_0/ca
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/array_obj_ref_1108_Merge/$entry
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/array_obj_ref_1108_Merge/$exit
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/array_obj_ref_1108_Merge/merge_req
      -- CP-element group 119: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1108_Update/array_obj_ref_1108_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1108_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1108_load_0_ack_1, ack => mainAcc2_CP_4584_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	0 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_sample_completed_
      -- CP-element group 120: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/$exit
      -- CP-element group 120: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/$exit
      -- CP-element group 120: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1111_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1111_load_0_ack_0, ack => mainAcc2_CP_4584_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	0 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	115 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_update_completed_
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/$exit
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/$exit
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/$entry
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/$exit
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/merge_req
      -- CP-element group 121: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1111_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1111_load_0_ack_1, ack => mainAcc2_CP_4584_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_sample_completed_
      -- CP-element group 122: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1113_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1113_inst_ack_0, ack => mainAcc2_CP_4584_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	0 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	151 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_update_completed_
      -- CP-element group 123: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Update/$exit
      -- CP-element group 123: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1113_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1113_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1113_inst_ack_1, ack => mainAcc2_CP_4584_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	130 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_sample_start_
      -- CP-element group 124: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1123_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(124), ack => type_cast_1123_inst_req_0); -- 
    mainAcc2_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(128) & mainAcc2_CP_4584_elements(130);
      gj_mainAcc2_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	6 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	196 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1118_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	0 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (18) 
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_sample_start_
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_word_address_calculated
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_root_address_calculated
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_offset_calculated
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_base_plus_offset/$entry
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_base_plus_offset/$exit
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_word_addrgen/$entry
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_word_addrgen/$exit
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_word_addrgen/root_register_req
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_word_addrgen/root_register_ack
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/$entry
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/$entry
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1118_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(126)); -- 
    rr_6222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(126), ack => array_obj_ref_1118_load_0_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_sample_completed_
      -- CP-element group 127: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/$exit
      -- CP-element group 127: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/$exit
      -- CP-element group 127: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/word_0/$exit
      -- CP-element group 127: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1118_load_0_ack_0, ack => mainAcc2_CP_4584_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	0 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	124 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_update_completed_
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/$exit
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/$exit
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/word_0/$exit
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/word_access_complete/word_0/ca
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/array_obj_ref_1118_Merge/$entry
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/array_obj_ref_1118_Merge/$exit
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/array_obj_ref_1118_Merge/merge_req
      -- CP-element group 128: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1118_Update/array_obj_ref_1118_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1118_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1118_load_0_ack_1, ack => mainAcc2_CP_4584_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	0 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_sample_completed_
      -- CP-element group 129: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/$exit
      -- CP-element group 129: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/$exit
      -- CP-element group 129: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/word_0/$exit
      -- CP-element group 129: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(129) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1121_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1121_load_0_ack_0, ack => mainAcc2_CP_4584_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	0 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	124 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_update_completed_
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/$exit
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/$exit
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/word_0/$exit
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/word_access_complete/word_0/ca
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/array_obj_ref_1121_Merge/$entry
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/array_obj_ref_1121_Merge/$exit
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/array_obj_ref_1121_Merge/merge_req
      -- CP-element group 130: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1121_Update/array_obj_ref_1121_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(130) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1121_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1121_load_0_ack_1, ack => mainAcc2_CP_4584_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	124 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_sample_completed_
      -- CP-element group 131: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Sample/$exit
      -- CP-element group 131: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(131) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1123_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_0, ack => mainAcc2_CP_4584_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	0 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	157 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_update_completed_
      -- CP-element group 132: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Update/$exit
      -- CP-element group 132: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1123_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(132) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1123_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1123_inst_ack_1, ack => mainAcc2_CP_4584_elements(132)); -- 
    -- CP-element group 133:  join  transition  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	139 
    -- CP-element group 133: 	137 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	140 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_sample_start_
      -- CP-element group 133: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Sample/$entry
      -- CP-element group 133: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(133) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1133_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(133), ack => type_cast_1133_inst_req_0); -- 
    mainAcc2_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(139) & mainAcc2_CP_4584_elements(137);
      gj_mainAcc2_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	6 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	196 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_sample_complete
      -- CP-element group 134: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(134) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	0 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (18) 
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_sample_start_
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_word_address_calculated
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_root_address_calculated
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_offset_calculated
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Update/$exit
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_final_index_sum_regn_Update/ack
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_base_plus_offset/$entry
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_base_plus_offset/$exit
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_base_plus_offset/sum_rename_req
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_base_plus_offset/sum_rename_ack
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_word_addrgen/$entry
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_word_addrgen/$exit
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_word_addrgen/root_register_req
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_word_addrgen/root_register_ack
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/$entry
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/$entry
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/word_0/$entry
      -- CP-element group 135: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(135)); -- 
    rr_6340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(135), ack => array_obj_ref_1128_load_0_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (5) 
      -- CP-element group 136: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_sample_completed_
      -- CP-element group 136: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/$exit
      -- CP-element group 136: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/$exit
      -- CP-element group 136: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/word_0/$exit
      -- CP-element group 136: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_load_0_ack_0, ack => mainAcc2_CP_4584_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	0 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (9) 
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_update_completed_
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/$exit
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/$exit
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/word_0/$exit
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/word_access_complete/word_0/ca
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/array_obj_ref_1128_Merge/$entry
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/array_obj_ref_1128_Merge/$exit
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/array_obj_ref_1128_Merge/merge_req
      -- CP-element group 137: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1128_Update/array_obj_ref_1128_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(137) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1128_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_load_0_ack_1, ack => mainAcc2_CP_4584_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	0 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (5) 
      -- CP-element group 138: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_sample_completed_
      -- CP-element group 138: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/$exit
      -- CP-element group 138: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/word_0/$exit
      -- CP-element group 138: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(138)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(138)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(138) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1131_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1131_load_0_ack_0, ack => mainAcc2_CP_4584_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	0 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	133 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_update_completed_
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/$exit
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/$exit
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/word_0/$exit
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/word_access_complete/word_0/ca
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/array_obj_ref_1131_Merge/$entry
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/array_obj_ref_1131_Merge/$exit
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/array_obj_ref_1131_Merge/merge_req
      -- CP-element group 139: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1131_Update/array_obj_ref_1131_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(139)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(139)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(139) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1131_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1131_load_0_ack_1, ack => mainAcc2_CP_4584_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	133 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_sample_completed_
      -- CP-element group 140: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Sample/$exit
      -- CP-element group 140: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(140)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(140)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(140) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1133_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1133_inst_ack_0, ack => mainAcc2_CP_4584_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	0 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	163 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_update_completed_
      -- CP-element group 141: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Update/$exit
      -- CP-element group 141: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1133_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(141)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(141)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(141) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1133_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1133_inst_ack_1, ack => mainAcc2_CP_4584_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	146 
    -- CP-element group 142: 	148 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	149 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_sample_start_
      -- CP-element group 142: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Sample/$entry
      -- CP-element group 142: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(142)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(142)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(142) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1143_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(142), ack => type_cast_1143_inst_req_0); -- 
    mainAcc2_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(146) & mainAcc2_CP_4584_elements(148);
      gj_mainAcc2_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	6 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	196 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_sample_complete
      -- CP-element group 143: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Sample/$exit
      -- CP-element group 143: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Sample/ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(143)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(143)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(143) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_index_offset_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1138_index_offset_ack_0, ack => mainAcc2_CP_4584_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	0 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (18) 
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_sample_start_
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_word_address_calculated
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_root_address_calculated
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_offset_calculated
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Update/$exit
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_final_index_sum_regn_Update/ack
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_base_plus_offset/$entry
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_base_plus_offset/$exit
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_base_plus_offset/sum_rename_req
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_base_plus_offset/sum_rename_ack
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_word_addrgen/$entry
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_word_addrgen/$exit
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_word_addrgen/root_register_req
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_word_addrgen/root_register_ack
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/$entry
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/$entry
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/word_0/$entry
      -- CP-element group 144: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(144)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(144)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(144) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_index_offset_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_6438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1138_index_offset_ack_1, ack => mainAcc2_CP_4584_elements(144)); -- 
    rr_6458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(144), ack => array_obj_ref_1138_load_0_req_0); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_sample_completed_
      -- CP-element group 145: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/$exit
      -- CP-element group 145: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/$exit
      -- CP-element group 145: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(145)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(145)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(145) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1138_load_0_ack_0, ack => mainAcc2_CP_4584_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	0 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	142 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_update_completed_
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/$exit
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/$exit
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/array_obj_ref_1138_Merge/$entry
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/array_obj_ref_1138_Merge/$exit
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/array_obj_ref_1138_Merge/merge_req
      -- CP-element group 146: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1138_Update/array_obj_ref_1138_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(146)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(146)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(146) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1138_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1138_load_0_ack_1, ack => mainAcc2_CP_4584_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	0 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_sample_completed_
      -- CP-element group 147: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/$exit
      -- CP-element group 147: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/$exit
      -- CP-element group 147: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/word_0/$exit
      -- CP-element group 147: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(147)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(147)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(147) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1141_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1141_load_0_ack_0, ack => mainAcc2_CP_4584_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	0 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	142 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_update_completed_
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/$exit
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/$exit
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/word_0/$exit
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/word_access_complete/word_0/ca
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/array_obj_ref_1141_Merge/$entry
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/array_obj_ref_1141_Merge/$exit
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/array_obj_ref_1141_Merge/merge_req
      -- CP-element group 148: 	 assign_stmt_934_to_assign_stmt_1234/array_obj_ref_1141_Update/array_obj_ref_1141_Merge/merge_ack
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(148)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(148)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(148) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:array_obj_ref_1141_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1141_load_0_ack_1, ack => mainAcc2_CP_4584_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	142 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_sample_completed_
      -- CP-element group 149: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Sample/$exit
      -- CP-element group 149: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(149)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(149)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(149) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1143_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1143_inst_ack_0, ack => mainAcc2_CP_4584_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	0 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	169 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_update_completed_
      -- CP-element group 150: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Update/$exit
      -- CP-element group 150: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1143_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(150)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(150)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(150) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1143_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1143_inst_ack_1, ack => mainAcc2_CP_4584_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	87 
    -- CP-element group 151: 	123 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_sample_start_
      -- CP-element group 151: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Sample/$entry
      -- CP-element group 151: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(151)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(151)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(151) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1149_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(151), ack => type_cast_1149_inst_req_0); -- 
    mainAcc2_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(87) & mainAcc2_CP_4584_elements(123);
      gj_mainAcc2_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_sample_completed_
      -- CP-element group 152: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Sample/$exit
      -- CP-element group 152: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(152)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(152)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(152) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1149_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_0, ack => mainAcc2_CP_4584_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	0 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	175 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_update_completed_
      -- CP-element group 153: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Update/$exit
      -- CP-element group 153: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1149_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(153)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(153)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(153) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1149_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_1, ack => mainAcc2_CP_4584_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	15 
    -- CP-element group 154: 	51 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_sample_start_
      -- CP-element group 154: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Sample/$entry
      -- CP-element group 154: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(154)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(154)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(154) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1155_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(154), ack => type_cast_1155_inst_req_0); -- 
    mainAcc2_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(15) & mainAcc2_CP_4584_elements(51);
      gj_mainAcc2_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_sample_completed_
      -- CP-element group 155: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Sample/$exit
      -- CP-element group 155: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(155)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(155)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(155) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1155_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_0, ack => mainAcc2_CP_4584_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	0 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	175 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_update_completed_
      -- CP-element group 156: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Update/$exit
      -- CP-element group 156: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1155_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(156)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(156)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(156) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1155_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1155_inst_ack_1, ack => mainAcc2_CP_4584_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	96 
    -- CP-element group 157: 	132 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_sample_start_
      -- CP-element group 157: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Sample/$entry
      -- CP-element group 157: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(157)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(157)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(157) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1161_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(157), ack => type_cast_1161_inst_req_0); -- 
    mainAcc2_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(96) & mainAcc2_CP_4584_elements(132);
      gj_mainAcc2_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_sample_completed_
      -- CP-element group 158: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Sample/$exit
      -- CP-element group 158: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(158)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(158)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(158) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1161_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_0, ack => mainAcc2_CP_4584_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	0 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	178 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_update_completed_
      -- CP-element group 159: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Update/$exit
      -- CP-element group 159: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1161_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(159)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(159)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(159) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1161_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_1, ack => mainAcc2_CP_4584_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	60 
    -- CP-element group 160: 	24 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_sample_start_
      -- CP-element group 160: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(160)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(160)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(160) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1167_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(160), ack => type_cast_1167_inst_req_0); -- 
    mainAcc2_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(60) & mainAcc2_CP_4584_elements(24);
      gj_mainAcc2_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_sample_completed_
      -- CP-element group 161: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Sample/$exit
      -- CP-element group 161: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(161)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(161)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(161) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1167_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => mainAcc2_CP_4584_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	0 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	178 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_update_completed_
      -- CP-element group 162: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Update/$exit
      -- CP-element group 162: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1167_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(162)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(162)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(162) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1167_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => mainAcc2_CP_4584_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	105 
    -- CP-element group 163: 	141 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_sample_start_
      -- CP-element group 163: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Sample/$entry
      -- CP-element group 163: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(163)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(163)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(163) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1173_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(163), ack => type_cast_1173_inst_req_0); -- 
    mainAcc2_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(105) & mainAcc2_CP_4584_elements(141);
      gj_mainAcc2_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_sample_completed_
      -- CP-element group 164: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Sample/$exit
      -- CP-element group 164: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(164)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(164)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(164) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1173_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => mainAcc2_CP_4584_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	0 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	181 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_update_completed_
      -- CP-element group 165: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Update/$exit
      -- CP-element group 165: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1173_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(165)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(165)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(165) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1173_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => mainAcc2_CP_4584_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	69 
    -- CP-element group 166: 	33 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_sample_start_
      -- CP-element group 166: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Sample/$entry
      -- CP-element group 166: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(166)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(166)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(166) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1179_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(166), ack => type_cast_1179_inst_req_0); -- 
    mainAcc2_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(69) & mainAcc2_CP_4584_elements(33);
      gj_mainAcc2_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_sample_completed_
      -- CP-element group 167: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Sample/$exit
      -- CP-element group 167: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(167)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(167)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(167) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1179_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_0, ack => mainAcc2_CP_4584_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	0 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	181 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_update_completed_
      -- CP-element group 168: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Update/$exit
      -- CP-element group 168: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1179_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(168)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(168)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(168) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1179_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_1, ack => mainAcc2_CP_4584_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	150 
    -- CP-element group 169: 	114 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_sample_start_
      -- CP-element group 169: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Sample/$entry
      -- CP-element group 169: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(169)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(169)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(169) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1185_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(169), ack => type_cast_1185_inst_req_0); -- 
    mainAcc2_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(150) & mainAcc2_CP_4584_elements(114);
      gj_mainAcc2_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_sample_completed_
      -- CP-element group 170: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Sample/$exit
      -- CP-element group 170: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(170)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(170)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(170) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1185_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1185_inst_ack_0, ack => mainAcc2_CP_4584_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	0 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	184 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_update_completed_
      -- CP-element group 171: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Update/$exit
      -- CP-element group 171: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1185_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(171)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(171)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(171) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1185_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1185_inst_ack_1, ack => mainAcc2_CP_4584_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	78 
    -- CP-element group 172: 	42 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_sample_start_
      -- CP-element group 172: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(172)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(172)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(172) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1191_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(172), ack => type_cast_1191_inst_req_0); -- 
    mainAcc2_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(78) & mainAcc2_CP_4584_elements(42);
      gj_mainAcc2_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_sample_completed_
      -- CP-element group 173: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Sample/$exit
      -- CP-element group 173: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(173)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(173)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(173) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1191_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_0, ack => mainAcc2_CP_4584_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	0 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	184 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_update_completed_
      -- CP-element group 174: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Update/$exit
      -- CP-element group 174: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1191_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(174)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(174)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(174) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1191_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1191_inst_ack_1, ack => mainAcc2_CP_4584_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	156 
    -- CP-element group 175: 	153 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_sample_start_
      -- CP-element group 175: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Sample/$entry
      -- CP-element group 175: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(175)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(175)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(175) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1197_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(175), ack => type_cast_1197_inst_req_0); -- 
    mainAcc2_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(156) & mainAcc2_CP_4584_elements(153);
      gj_mainAcc2_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_sample_completed_
      -- CP-element group 176: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Sample/$exit
      -- CP-element group 176: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(176)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(176)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(176) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1197_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_0, ack => mainAcc2_CP_4584_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	0 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	187 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_update_completed_
      -- CP-element group 177: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Update/$exit
      -- CP-element group 177: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1197_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(177)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(177)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(177) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1197_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_1, ack => mainAcc2_CP_4584_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	162 
    -- CP-element group 178: 	159 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_sample_start_
      -- CP-element group 178: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Sample/$entry
      -- CP-element group 178: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(178)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(178)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(178) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1203_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(178), ack => type_cast_1203_inst_req_0); -- 
    mainAcc2_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(162) & mainAcc2_CP_4584_elements(159);
      gj_mainAcc2_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_sample_completed_
      -- CP-element group 179: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Sample/$exit
      -- CP-element group 179: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(179)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(179)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(179) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1203_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_0, ack => mainAcc2_CP_4584_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	0 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	187 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_update_completed_
      -- CP-element group 180: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Update/$exit
      -- CP-element group 180: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1203_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(180)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(180)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(180) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1203_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_1, ack => mainAcc2_CP_4584_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	168 
    -- CP-element group 181: 	165 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_sample_start_
      -- CP-element group 181: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Sample/$entry
      -- CP-element group 181: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(181)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(181)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(181) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1209_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(181), ack => type_cast_1209_inst_req_0); -- 
    mainAcc2_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(168) & mainAcc2_CP_4584_elements(165);
      gj_mainAcc2_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_sample_completed_
      -- CP-element group 182: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Sample/$exit
      -- CP-element group 182: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(182)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(182)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(182) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1209_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_0, ack => mainAcc2_CP_4584_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	0 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	190 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_update_completed_
      -- CP-element group 183: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Update/$exit
      -- CP-element group 183: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1209_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(183)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(183)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(183) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1209_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_1, ack => mainAcc2_CP_4584_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	171 
    -- CP-element group 184: 	174 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_sample_start_
      -- CP-element group 184: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Sample/$entry
      -- CP-element group 184: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(184)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(184)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(184) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1215_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(184), ack => type_cast_1215_inst_req_0); -- 
    mainAcc2_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(171) & mainAcc2_CP_4584_elements(174);
      gj_mainAcc2_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_sample_completed_
      -- CP-element group 185: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Sample/$exit
      -- CP-element group 185: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(185)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(185)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(185) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1215_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_0, ack => mainAcc2_CP_4584_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	0 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	190 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_update_completed_
      -- CP-element group 186: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Update/$exit
      -- CP-element group 186: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1215_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(186)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(186)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(186) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1215_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1215_inst_ack_1, ack => mainAcc2_CP_4584_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	180 
    -- CP-element group 187: 	177 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_sample_start_
      -- CP-element group 187: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Sample/$entry
      -- CP-element group 187: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(187)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(187)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(187) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1221_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(187), ack => type_cast_1221_inst_req_0); -- 
    mainAcc2_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(180) & mainAcc2_CP_4584_elements(177);
      gj_mainAcc2_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_sample_completed_
      -- CP-element group 188: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Sample/$exit
      -- CP-element group 188: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(188)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(188)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(188) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1221_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => mainAcc2_CP_4584_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	0 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	193 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_update_completed_
      -- CP-element group 189: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Update/$exit
      -- CP-element group 189: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1221_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(189)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(189)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(189) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1221_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => mainAcc2_CP_4584_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	186 
    -- CP-element group 190: 	183 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_sample_start_
      -- CP-element group 190: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Sample/$entry
      -- CP-element group 190: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(190)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(190)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(190) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1227_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(190), ack => type_cast_1227_inst_req_0); -- 
    mainAcc2_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(186) & mainAcc2_CP_4584_elements(183);
      gj_mainAcc2_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_sample_completed_
      -- CP-element group 191: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Sample/$exit
      -- CP-element group 191: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(191)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(191)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(191) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1227_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_0, ack => mainAcc2_CP_4584_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	0 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_update_completed_
      -- CP-element group 192: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Update/$exit
      -- CP-element group 192: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1227_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(192)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(192)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(192) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1227_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1227_inst_ack_1, ack => mainAcc2_CP_4584_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	189 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_sample_start_
      -- CP-element group 193: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Sample/$entry
      -- CP-element group 193: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Sample/rr
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(193)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(193)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(193) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1233_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_6723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => mainAcc2_CP_4584_elements(193), ack => type_cast_1233_inst_req_0); -- 
    mainAcc2_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(192) & mainAcc2_CP_4584_elements(189);
      gj_mainAcc2_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_sample_completed_
      -- CP-element group 194: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Sample/ra
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(194)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(194)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(194) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1233_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_6724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_0, ack => mainAcc2_CP_4584_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	0 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_update_completed_
      -- CP-element group 195: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Update/$exit
      -- CP-element group 195: 	 assign_stmt_934_to_assign_stmt_1234/type_cast_1233_Update/ca
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(195)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(195)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(195) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:type_cast_1233_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_6729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1233_inst_ack_1, ack => mainAcc2_CP_4584_elements(195)); -- 
    -- CP-element group 196:  join  transition  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	89 
    -- CP-element group 196: 	44 
    -- CP-element group 196: 	53 
    -- CP-element group 196: 	26 
    -- CP-element group 196: 	62 
    -- CP-element group 196: 	8 
    -- CP-element group 196: 	17 
    -- CP-element group 196: 	71 
    -- CP-element group 196: 	80 
    -- CP-element group 196: 	98 
    -- CP-element group 196: 	107 
    -- CP-element group 196: 	195 
    -- CP-element group 196: 	35 
    -- CP-element group 196: 	143 
    -- CP-element group 196: 	125 
    -- CP-element group 196: 	134 
    -- CP-element group 196: 	116 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 $exit
      -- CP-element group 196: 	 assign_stmt_934_to_assign_stmt_1234/$exit
      -- 
    -- logger for CP element group mainAcc2_CP_4584_elements(196)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and mainAcc2_CP_4584_elements(196)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:mainAcc2:CP:mainAcc2_CP_4584_elements(196) fired."); 
        -- 
      end if; --
    end process; 
    mainAcc2_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 29) := "mainAcc2_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= mainAcc2_CP_4584_elements(89) & mainAcc2_CP_4584_elements(44) & mainAcc2_CP_4584_elements(53) & mainAcc2_CP_4584_elements(26) & mainAcc2_CP_4584_elements(62) & mainAcc2_CP_4584_elements(8) & mainAcc2_CP_4584_elements(17) & mainAcc2_CP_4584_elements(71) & mainAcc2_CP_4584_elements(80) & mainAcc2_CP_4584_elements(98) & mainAcc2_CP_4584_elements(107) & mainAcc2_CP_4584_elements(195) & mainAcc2_CP_4584_elements(35) & mainAcc2_CP_4584_elements(143) & mainAcc2_CP_4584_elements(125) & mainAcc2_CP_4584_elements(134) & mainAcc2_CP_4584_elements(116);
      gj_mainAcc2_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => mainAcc2_CP_4584_elements(196), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1148_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1154_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1160_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1166_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1172_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1178_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1184_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1190_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1196_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1202_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1208_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1214_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1220_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1226_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_1232_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_969_wire : std_logic_vector(1 downto 0);
    signal ADD_u2_u2_981_wire : std_logic_vector(1 downto 0);
    signal EQ_u2_u1_950_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_976_wire : std_logic_vector(0 downto 0);
    signal MUL_u16_u16_1002_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1012_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1022_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1032_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1042_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1052_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1062_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1072_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1082_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1092_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1102_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1112_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1122_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1132_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_1142_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_992_wire : std_logic_vector(15 downto 0);
    signal R_col_to_be_replaced_1007_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1007_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1017_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1017_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1027_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1027_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1037_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1037_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1047_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1047_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1057_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_1_1057_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1067_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1067_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1077_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1077_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1087_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1087_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1097_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_2_1097_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1107_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1107_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1117_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1117_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1127_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1127_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1137_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_3_1137_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_987_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_987_scaled : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_997_resized : std_logic_vector(3 downto 0);
    signal R_col_to_be_replaced_997_scaled : std_logic_vector(3 downto 0);
    signal SUB_u2_u2_955_wire : std_logic_vector(1 downto 0);
    signal SUB_u2_u2_965_wire : std_logic_vector(1 downto 0);
    signal UGE_u2_u1_962_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_1001_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1001_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1001_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1008_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1008_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1008_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1011_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1011_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1011_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1018_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1018_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1018_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1021_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1021_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1021_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1028_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1028_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1028_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1031_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1031_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1031_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1038_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1038_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1038_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1041_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1041_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1041_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1048_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1051_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1051_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1051_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1058_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1058_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1058_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1061_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1061_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1061_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1068_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1068_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1068_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1071_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1071_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1071_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1078_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1078_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1078_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1081_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1081_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1081_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1088_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1088_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1088_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1091_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1091_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1091_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1098_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1098_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1098_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1101_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1101_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1101_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1108_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1108_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1108_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1111_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1111_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1111_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1118_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1118_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1118_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1121_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1121_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1121_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1128_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1128_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1128_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1131_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1131_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1131_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1138_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1138_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1138_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_1141_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1141_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_1141_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_988_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_988_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_988_word_offset_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_991_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_991_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_991_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_constant_part_of_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_data_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_998_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_offset_scale_factor_1 : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_wire : std_logic_vector(15 downto 0);
    signal array_obj_ref_998_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_998_word_offset_0 : std_logic_vector(3 downto 0);
    signal col_to_be_replaced_1_958 : std_logic_vector(1 downto 0);
    signal col_to_be_replaced_2_972 : std_logic_vector(1 downto 0);
    signal col_to_be_replaced_3_984 : std_logic_vector(1 downto 0);
    signal konst_949_wire_constant : std_logic_vector(1 downto 0);
    signal konst_954_wire_constant : std_logic_vector(1 downto 0);
    signal konst_961_wire_constant : std_logic_vector(1 downto 0);
    signal konst_964_wire_constant : std_logic_vector(1 downto 0);
    signal konst_968_wire_constant : std_logic_vector(1 downto 0);
    signal konst_975_wire_constant : std_logic_vector(1 downto 0);
    signal konst_980_wire_constant : std_logic_vector(1 downto 0);
    signal one_938 : std_logic_vector(1 downto 0);
    signal pp00_1114 : std_logic_vector(15 downto 0);
    signal pp01_1074 : std_logic_vector(15 downto 0);
    signal pp02_1034 : std_logic_vector(15 downto 0);
    signal pp03_994 : std_logic_vector(15 downto 0);
    signal pp10_1124 : std_logic_vector(15 downto 0);
    signal pp11_1084 : std_logic_vector(15 downto 0);
    signal pp12_1044 : std_logic_vector(15 downto 0);
    signal pp13_1004 : std_logic_vector(15 downto 0);
    signal pp20_1134 : std_logic_vector(15 downto 0);
    signal pp21_1094 : std_logic_vector(15 downto 0);
    signal pp22_1054 : std_logic_vector(15 downto 0);
    signal pp23_1014 : std_logic_vector(15 downto 0);
    signal pp30_1144 : std_logic_vector(15 downto 0);
    signal pp31_1104 : std_logic_vector(15 downto 0);
    signal pp32_1064 : std_logic_vector(15 downto 0);
    signal pp33_1024 : std_logic_vector(15 downto 0);
    signal sum0_1150 : std_logic_vector(15 downto 0);
    signal sum10_1198 : std_logic_vector(15 downto 0);
    signal sum11_1204 : std_logic_vector(15 downto 0);
    signal sum12_1210 : std_logic_vector(15 downto 0);
    signal sum13_1216 : std_logic_vector(15 downto 0);
    signal sum1_1156 : std_logic_vector(15 downto 0);
    signal sum20_1222 : std_logic_vector(15 downto 0);
    signal sum21_1228 : std_logic_vector(15 downto 0);
    signal sum2_1162 : std_logic_vector(15 downto 0);
    signal sum3_1168 : std_logic_vector(15 downto 0);
    signal sum4_1174 : std_logic_vector(15 downto 0);
    signal sum5_1180 : std_logic_vector(15 downto 0);
    signal sum6_1186 : std_logic_vector(15 downto 0);
    signal sum7_1192 : std_logic_vector(15 downto 0);
    signal three_946 : std_logic_vector(1 downto 0);
    signal two_942 : std_logic_vector(1 downto 0);
    signal type_cast_952_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_956_wire : std_logic_vector(1 downto 0);
    signal type_cast_966_wire : std_logic_vector(1 downto 0);
    signal type_cast_970_wire : std_logic_vector(1 downto 0);
    signal type_cast_978_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_982_wire : std_logic_vector(1 downto 0);
    signal zero_934 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_1001_word_address_0 <= "0111";
    array_obj_ref_1008_constant_part_of_offset <= "1000";
    array_obj_ref_1008_offset_scale_factor_0 <= "0100";
    array_obj_ref_1008_offset_scale_factor_1 <= "0001";
    array_obj_ref_1008_resized_base_address <= "0000";
    array_obj_ref_1008_word_offset_0 <= "0000";
    array_obj_ref_1011_word_address_0 <= "1011";
    array_obj_ref_1018_constant_part_of_offset <= "1100";
    array_obj_ref_1018_offset_scale_factor_0 <= "0100";
    array_obj_ref_1018_offset_scale_factor_1 <= "0001";
    array_obj_ref_1018_resized_base_address <= "0000";
    array_obj_ref_1018_word_offset_0 <= "0000";
    array_obj_ref_1021_word_address_0 <= "1111";
    array_obj_ref_1028_constant_part_of_offset <= "0000";
    array_obj_ref_1028_offset_scale_factor_0 <= "0100";
    array_obj_ref_1028_offset_scale_factor_1 <= "0001";
    array_obj_ref_1028_resized_base_address <= "0000";
    array_obj_ref_1028_word_offset_0 <= "0000";
    array_obj_ref_1031_word_address_0 <= "0010";
    array_obj_ref_1038_constant_part_of_offset <= "0100";
    array_obj_ref_1038_offset_scale_factor_0 <= "0100";
    array_obj_ref_1038_offset_scale_factor_1 <= "0001";
    array_obj_ref_1038_resized_base_address <= "0000";
    array_obj_ref_1038_word_offset_0 <= "0000";
    array_obj_ref_1041_word_address_0 <= "0110";
    array_obj_ref_1048_constant_part_of_offset <= "1000";
    array_obj_ref_1048_offset_scale_factor_0 <= "0100";
    array_obj_ref_1048_offset_scale_factor_1 <= "0001";
    array_obj_ref_1048_resized_base_address <= "0000";
    array_obj_ref_1048_word_offset_0 <= "0000";
    array_obj_ref_1051_word_address_0 <= "1010";
    array_obj_ref_1058_constant_part_of_offset <= "1100";
    array_obj_ref_1058_offset_scale_factor_0 <= "0100";
    array_obj_ref_1058_offset_scale_factor_1 <= "0001";
    array_obj_ref_1058_resized_base_address <= "0000";
    array_obj_ref_1058_word_offset_0 <= "0000";
    array_obj_ref_1061_word_address_0 <= "1110";
    array_obj_ref_1068_constant_part_of_offset <= "0000";
    array_obj_ref_1068_offset_scale_factor_0 <= "0100";
    array_obj_ref_1068_offset_scale_factor_1 <= "0001";
    array_obj_ref_1068_resized_base_address <= "0000";
    array_obj_ref_1068_word_offset_0 <= "0000";
    array_obj_ref_1071_word_address_0 <= "0001";
    array_obj_ref_1078_constant_part_of_offset <= "0100";
    array_obj_ref_1078_offset_scale_factor_0 <= "0100";
    array_obj_ref_1078_offset_scale_factor_1 <= "0001";
    array_obj_ref_1078_resized_base_address <= "0000";
    array_obj_ref_1078_word_offset_0 <= "0000";
    array_obj_ref_1081_word_address_0 <= "0101";
    array_obj_ref_1088_constant_part_of_offset <= "1000";
    array_obj_ref_1088_offset_scale_factor_0 <= "0100";
    array_obj_ref_1088_offset_scale_factor_1 <= "0001";
    array_obj_ref_1088_resized_base_address <= "0000";
    array_obj_ref_1088_word_offset_0 <= "0000";
    array_obj_ref_1091_word_address_0 <= "1001";
    array_obj_ref_1098_constant_part_of_offset <= "1100";
    array_obj_ref_1098_offset_scale_factor_0 <= "0100";
    array_obj_ref_1098_offset_scale_factor_1 <= "0001";
    array_obj_ref_1098_resized_base_address <= "0000";
    array_obj_ref_1098_word_offset_0 <= "0000";
    array_obj_ref_1101_word_address_0 <= "1101";
    array_obj_ref_1108_constant_part_of_offset <= "0000";
    array_obj_ref_1108_offset_scale_factor_0 <= "0100";
    array_obj_ref_1108_offset_scale_factor_1 <= "0001";
    array_obj_ref_1108_resized_base_address <= "0000";
    array_obj_ref_1108_word_offset_0 <= "0000";
    array_obj_ref_1111_word_address_0 <= "0000";
    array_obj_ref_1118_constant_part_of_offset <= "0100";
    array_obj_ref_1118_offset_scale_factor_0 <= "0100";
    array_obj_ref_1118_offset_scale_factor_1 <= "0001";
    array_obj_ref_1118_resized_base_address <= "0000";
    array_obj_ref_1118_word_offset_0 <= "0000";
    array_obj_ref_1121_word_address_0 <= "0100";
    array_obj_ref_1128_constant_part_of_offset <= "1000";
    array_obj_ref_1128_offset_scale_factor_0 <= "0100";
    array_obj_ref_1128_offset_scale_factor_1 <= "0001";
    array_obj_ref_1128_resized_base_address <= "0000";
    array_obj_ref_1128_word_offset_0 <= "0000";
    array_obj_ref_1131_word_address_0 <= "1000";
    array_obj_ref_1138_constant_part_of_offset <= "1100";
    array_obj_ref_1138_offset_scale_factor_0 <= "0100";
    array_obj_ref_1138_offset_scale_factor_1 <= "0001";
    array_obj_ref_1138_resized_base_address <= "0000";
    array_obj_ref_1138_word_offset_0 <= "0000";
    array_obj_ref_1141_word_address_0 <= "1100";
    array_obj_ref_988_constant_part_of_offset <= "0000";
    array_obj_ref_988_offset_scale_factor_0 <= "0100";
    array_obj_ref_988_offset_scale_factor_1 <= "0001";
    array_obj_ref_988_resized_base_address <= "0000";
    array_obj_ref_988_word_offset_0 <= "0000";
    array_obj_ref_991_word_address_0 <= "0011";
    array_obj_ref_998_constant_part_of_offset <= "0100";
    array_obj_ref_998_offset_scale_factor_0 <= "0100";
    array_obj_ref_998_offset_scale_factor_1 <= "0001";
    array_obj_ref_998_resized_base_address <= "0000";
    array_obj_ref_998_word_offset_0 <= "0000";
    konst_949_wire_constant <= "00";
    konst_954_wire_constant <= "01";
    konst_961_wire_constant <= "10";
    konst_964_wire_constant <= "10";
    konst_968_wire_constant <= "10";
    konst_975_wire_constant <= "11";
    konst_980_wire_constant <= "01";
    one_938 <= "01";
    three_946 <= "11";
    two_942 <= "10";
    type_cast_952_wire_constant <= "11";
    type_cast_978_wire_constant <= "00";
    zero_934 <= "00";
    -- logger for split-operator MUX_957_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_957_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_957_inst:started:   inputs: " & " EQ_u2_u1_950_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_950_wire) & " type_cast_952_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_952_wire_constant) & " type_cast_956_wire = "& Convert_SLV_To_Hex_String(type_cast_956_wire));
          --
        end if; 
        if MUX_957_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_957_inst:finished:  outputs: " & " col_to_be_replaced_1_958= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_1_958));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_957_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_957_inst_req_0;
      MUX_957_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_957_inst_req_1;
      MUX_957_inst_ack_1<= update_ack(0);
      MUX_957_inst: SelectSplitProtocol generic map(name => "MUX_957_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_952_wire_constant, y => type_cast_956_wire, sel => EQ_u2_u1_950_wire, z => col_to_be_replaced_1_958, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_971_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_971_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_971_inst:started:   inputs: " & " UGE_u2_u1_962_wire = "& Convert_SLV_To_Hex_String(UGE_u2_u1_962_wire) & " type_cast_966_wire = "& Convert_SLV_To_Hex_String(type_cast_966_wire) & " type_cast_970_wire = "& Convert_SLV_To_Hex_String(type_cast_970_wire));
          --
        end if; 
        if MUX_971_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_971_inst:finished:  outputs: " & " col_to_be_replaced_2_972= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_2_972));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_971_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_971_inst_req_0;
      MUX_971_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_971_inst_req_1;
      MUX_971_inst_ack_1<= update_ack(0);
      MUX_971_inst: SelectSplitProtocol generic map(name => "MUX_971_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_966_wire, y => type_cast_970_wire, sel => UGE_u2_u1_962_wire, z => col_to_be_replaced_2_972, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator MUX_983_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_983_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_983_inst:started:   inputs: " & " EQ_u2_u1_976_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_976_wire) & " type_cast_978_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_978_wire_constant) & " type_cast_982_wire = "& Convert_SLV_To_Hex_String(type_cast_982_wire));
          --
        end if; 
        if MUX_983_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUX_983_inst:finished:  outputs: " & " col_to_be_replaced_3_984= "  & Convert_SLV_To_Hex_String(col_to_be_replaced_3_984));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_983_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_983_inst_req_0;
      MUX_983_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_983_inst_req_1;
      MUX_983_inst_ack_1<= update_ack(0);
      MUX_983_inst: SelectSplitProtocol generic map(name => "MUX_983_inst", data_width => 2, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => type_cast_978_wire_constant, y => type_cast_982_wire, sel => EQ_u2_u1_976_wire, z => col_to_be_replaced_3_984, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator type_cast_1003_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1003_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1003_inst:started:   inputs: " & " MUL_u16_u16_1002_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1002_wire));
          --
        end if; 
        if type_cast_1003_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1003_inst:finished:  outputs: " & " pp13_1004= "  & Convert_SLV_To_Hex_String(pp13_1004));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1003_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1003_inst_req_0;
      type_cast_1003_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1003_inst_req_1;
      type_cast_1003_inst_ack_1<= rack(0);
      type_cast_1003_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1003_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1002_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp13_1004,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1013_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1013_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1013_inst:started:   inputs: " & " MUL_u16_u16_1012_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1012_wire));
          --
        end if; 
        if type_cast_1013_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1013_inst:finished:  outputs: " & " pp23_1014= "  & Convert_SLV_To_Hex_String(pp23_1014));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1013_inst_req_0;
      type_cast_1013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1013_inst_req_1;
      type_cast_1013_inst_ack_1<= rack(0);
      type_cast_1013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1012_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp23_1014,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1023_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1023_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1023_inst:started:   inputs: " & " MUL_u16_u16_1022_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1022_wire));
          --
        end if; 
        if type_cast_1023_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1023_inst:finished:  outputs: " & " pp33_1024= "  & Convert_SLV_To_Hex_String(pp33_1024));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1023_inst_req_0;
      type_cast_1023_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1023_inst_req_1;
      type_cast_1023_inst_ack_1<= rack(0);
      type_cast_1023_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1023_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1022_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp33_1024,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1033_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1033_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1033_inst:started:   inputs: " & " MUL_u16_u16_1032_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1032_wire));
          --
        end if; 
        if type_cast_1033_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1033_inst:finished:  outputs: " & " pp02_1034= "  & Convert_SLV_To_Hex_String(pp02_1034));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1033_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1033_inst_req_0;
      type_cast_1033_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1033_inst_req_1;
      type_cast_1033_inst_ack_1<= rack(0);
      type_cast_1033_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1033_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1032_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp02_1034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1043_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1043_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1043_inst:started:   inputs: " & " MUL_u16_u16_1042_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1042_wire));
          --
        end if; 
        if type_cast_1043_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1043_inst:finished:  outputs: " & " pp12_1044= "  & Convert_SLV_To_Hex_String(pp12_1044));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1043_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1043_inst_req_0;
      type_cast_1043_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1043_inst_req_1;
      type_cast_1043_inst_ack_1<= rack(0);
      type_cast_1043_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1043_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1042_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp12_1044,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1053_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1053_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1053_inst:started:   inputs: " & " MUL_u16_u16_1052_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1052_wire));
          --
        end if; 
        if type_cast_1053_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1053_inst:finished:  outputs: " & " pp22_1054= "  & Convert_SLV_To_Hex_String(pp22_1054));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1053_inst_req_0;
      type_cast_1053_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1053_inst_req_1;
      type_cast_1053_inst_ack_1<= rack(0);
      type_cast_1053_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1053_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1052_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp22_1054,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1063_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1063_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1063_inst:started:   inputs: " & " MUL_u16_u16_1062_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1062_wire));
          --
        end if; 
        if type_cast_1063_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1063_inst:finished:  outputs: " & " pp32_1064= "  & Convert_SLV_To_Hex_String(pp32_1064));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1063_inst_req_0;
      type_cast_1063_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1063_inst_req_1;
      type_cast_1063_inst_ack_1<= rack(0);
      type_cast_1063_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1063_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1062_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp32_1064,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1073_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1073_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1073_inst:started:   inputs: " & " MUL_u16_u16_1072_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1072_wire));
          --
        end if; 
        if type_cast_1073_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1073_inst:finished:  outputs: " & " pp01_1074= "  & Convert_SLV_To_Hex_String(pp01_1074));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1073_inst_req_0;
      type_cast_1073_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1073_inst_req_1;
      type_cast_1073_inst_ack_1<= rack(0);
      type_cast_1073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1072_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp01_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1083_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1083_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1083_inst:started:   inputs: " & " MUL_u16_u16_1082_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1082_wire));
          --
        end if; 
        if type_cast_1083_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1083_inst:finished:  outputs: " & " pp11_1084= "  & Convert_SLV_To_Hex_String(pp11_1084));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1083_inst_req_0;
      type_cast_1083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1083_inst_req_1;
      type_cast_1083_inst_ack_1<= rack(0);
      type_cast_1083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1082_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp11_1084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1093_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1093_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1093_inst:started:   inputs: " & " MUL_u16_u16_1092_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1092_wire));
          --
        end if; 
        if type_cast_1093_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1093_inst:finished:  outputs: " & " pp21_1094= "  & Convert_SLV_To_Hex_String(pp21_1094));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1093_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1093_inst_req_0;
      type_cast_1093_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1093_inst_req_1;
      type_cast_1093_inst_ack_1<= rack(0);
      type_cast_1093_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1093_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1092_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp21_1094,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1103_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1103_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1103_inst:started:   inputs: " & " MUL_u16_u16_1102_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1102_wire));
          --
        end if; 
        if type_cast_1103_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1103_inst:finished:  outputs: " & " pp31_1104= "  & Convert_SLV_To_Hex_String(pp31_1104));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1103_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1103_inst_req_0;
      type_cast_1103_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1103_inst_req_1;
      type_cast_1103_inst_ack_1<= rack(0);
      type_cast_1103_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1103_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1102_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp31_1104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1113_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1113_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1113_inst:started:   inputs: " & " MUL_u16_u16_1112_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1112_wire));
          --
        end if; 
        if type_cast_1113_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1113_inst:finished:  outputs: " & " pp00_1114= "  & Convert_SLV_To_Hex_String(pp00_1114));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1113_inst_req_0;
      type_cast_1113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1113_inst_req_1;
      type_cast_1113_inst_ack_1<= rack(0);
      type_cast_1113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1112_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp00_1114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1123_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1123_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1123_inst:started:   inputs: " & " MUL_u16_u16_1122_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1122_wire));
          --
        end if; 
        if type_cast_1123_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1123_inst:finished:  outputs: " & " pp10_1124= "  & Convert_SLV_To_Hex_String(pp10_1124));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1123_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1123_inst_req_0;
      type_cast_1123_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1123_inst_req_1;
      type_cast_1123_inst_ack_1<= rack(0);
      type_cast_1123_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1123_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1122_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp10_1124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1133_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1133_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1133_inst:started:   inputs: " & " MUL_u16_u16_1132_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1132_wire));
          --
        end if; 
        if type_cast_1133_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1133_inst:finished:  outputs: " & " pp20_1134= "  & Convert_SLV_To_Hex_String(pp20_1134));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1133_inst_req_0;
      type_cast_1133_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1133_inst_req_1;
      type_cast_1133_inst_ack_1<= rack(0);
      type_cast_1133_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1133_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1132_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp20_1134,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1143_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1143_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1143_inst:started:   inputs: " & " MUL_u16_u16_1142_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_1142_wire));
          --
        end if; 
        if type_cast_1143_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1143_inst:finished:  outputs: " & " pp30_1144= "  & Convert_SLV_To_Hex_String(pp30_1144));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1143_inst_req_0;
      type_cast_1143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1143_inst_req_1;
      type_cast_1143_inst_ack_1<= rack(0);
      type_cast_1143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_1142_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp30_1144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1149_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1149_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1149_inst:started:   inputs: " & " ADD_u16_u16_1148_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1148_wire));
          --
        end if; 
        if type_cast_1149_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1149_inst:finished:  outputs: " & " sum0_1150= "  & Convert_SLV_To_Hex_String(sum0_1150));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1149_inst_req_0;
      type_cast_1149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1149_inst_req_1;
      type_cast_1149_inst_ack_1<= rack(0);
      type_cast_1149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1148_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum0_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1155_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1155_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1155_inst:started:   inputs: " & " ADD_u16_u16_1154_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1154_wire));
          --
        end if; 
        if type_cast_1155_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1155_inst:finished:  outputs: " & " sum1_1156= "  & Convert_SLV_To_Hex_String(sum1_1156));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1155_inst_req_0;
      type_cast_1155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1155_inst_req_1;
      type_cast_1155_inst_ack_1<= rack(0);
      type_cast_1155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1154_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum1_1156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1161_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1161_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1161_inst:started:   inputs: " & " ADD_u16_u16_1160_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1160_wire));
          --
        end if; 
        if type_cast_1161_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1161_inst:finished:  outputs: " & " sum2_1162= "  & Convert_SLV_To_Hex_String(sum2_1162));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1161_inst_req_0;
      type_cast_1161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1161_inst_req_1;
      type_cast_1161_inst_ack_1<= rack(0);
      type_cast_1161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1160_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum2_1162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1167_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1167_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1167_inst:started:   inputs: " & " ADD_u16_u16_1166_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1166_wire));
          --
        end if; 
        if type_cast_1167_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1167_inst:finished:  outputs: " & " sum3_1168= "  & Convert_SLV_To_Hex_String(sum3_1168));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1166_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum3_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1173_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1173_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1173_inst:started:   inputs: " & " ADD_u16_u16_1172_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1172_wire));
          --
        end if; 
        if type_cast_1173_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1173_inst:finished:  outputs: " & " sum4_1174= "  & Convert_SLV_To_Hex_String(sum4_1174));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1172_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum4_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1179_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1179_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1179_inst:started:   inputs: " & " ADD_u16_u16_1178_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1178_wire));
          --
        end if; 
        if type_cast_1179_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1179_inst:finished:  outputs: " & " sum5_1180= "  & Convert_SLV_To_Hex_String(sum5_1180));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1179_inst_req_0;
      type_cast_1179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1179_inst_req_1;
      type_cast_1179_inst_ack_1<= rack(0);
      type_cast_1179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1178_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum5_1180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1185_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1185_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1185_inst:started:   inputs: " & " ADD_u16_u16_1184_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1184_wire));
          --
        end if; 
        if type_cast_1185_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1185_inst:finished:  outputs: " & " sum6_1186= "  & Convert_SLV_To_Hex_String(sum6_1186));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1185_inst_req_0;
      type_cast_1185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1185_inst_req_1;
      type_cast_1185_inst_ack_1<= rack(0);
      type_cast_1185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1184_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum6_1186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1191_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1191_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1191_inst:started:   inputs: " & " ADD_u16_u16_1190_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1190_wire));
          --
        end if; 
        if type_cast_1191_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1191_inst:finished:  outputs: " & " sum7_1192= "  & Convert_SLV_To_Hex_String(sum7_1192));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1191_inst_req_0;
      type_cast_1191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1191_inst_req_1;
      type_cast_1191_inst_ack_1<= rack(0);
      type_cast_1191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1190_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum7_1192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1197_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1197_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1197_inst:started:   inputs: " & " ADD_u16_u16_1196_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1196_wire));
          --
        end if; 
        if type_cast_1197_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1197_inst:finished:  outputs: " & " sum10_1198= "  & Convert_SLV_To_Hex_String(sum10_1198));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1197_inst_req_0;
      type_cast_1197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1197_inst_req_1;
      type_cast_1197_inst_ack_1<= rack(0);
      type_cast_1197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1196_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum10_1198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1203_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1203_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1203_inst:started:   inputs: " & " ADD_u16_u16_1202_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1202_wire));
          --
        end if; 
        if type_cast_1203_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1203_inst:finished:  outputs: " & " sum11_1204= "  & Convert_SLV_To_Hex_String(sum11_1204));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1203_inst_req_0;
      type_cast_1203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1203_inst_req_1;
      type_cast_1203_inst_ack_1<= rack(0);
      type_cast_1203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1202_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum11_1204,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1209_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1209_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1209_inst:started:   inputs: " & " ADD_u16_u16_1208_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1208_wire));
          --
        end if; 
        if type_cast_1209_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1209_inst:finished:  outputs: " & " sum12_1210= "  & Convert_SLV_To_Hex_String(sum12_1210));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1209_inst_req_0;
      type_cast_1209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1209_inst_req_1;
      type_cast_1209_inst_ack_1<= rack(0);
      type_cast_1209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1208_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum12_1210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1215_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1215_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1215_inst:started:   inputs: " & " ADD_u16_u16_1214_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1214_wire));
          --
        end if; 
        if type_cast_1215_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1215_inst:finished:  outputs: " & " sum13_1216= "  & Convert_SLV_To_Hex_String(sum13_1216));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1215_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1215_inst_req_0;
      type_cast_1215_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1215_inst_req_1;
      type_cast_1215_inst_ack_1<= rack(0);
      type_cast_1215_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1215_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1214_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum13_1216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1221_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1221_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1221_inst:started:   inputs: " & " ADD_u16_u16_1220_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1220_wire));
          --
        end if; 
        if type_cast_1221_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1221_inst:finished:  outputs: " & " sum20_1222= "  & Convert_SLV_To_Hex_String(sum20_1222));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1220_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum20_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1227_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1227_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1227_inst:started:   inputs: " & " ADD_u16_u16_1226_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1226_wire));
          --
        end if; 
        if type_cast_1227_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1227_inst:finished:  outputs: " & " sum21_1228= "  & Convert_SLV_To_Hex_String(sum21_1228));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1227_inst_req_0;
      type_cast_1227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1227_inst_req_1;
      type_cast_1227_inst_ack_1<= rack(0);
      type_cast_1227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1226_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sum21_1228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1233_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1233_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1233_inst:started:   inputs: " & " ADD_u16_u16_1232_wire = "& Convert_SLV_To_Hex_String(ADD_u16_u16_1232_wire));
          --
        end if; 
        if type_cast_1233_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_1233_inst:finished:  outputs: " & " ofmap_pixel_buffer= "  & Convert_SLV_To_Hex_String(ofmap_pixel_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1233_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1233_inst_req_0;
      type_cast_1233_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1233_inst_req_1;
      type_cast_1233_inst_ack_1<= rack(0);
      type_cast_1233_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1233_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u16_u16_1232_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ofmap_pixel_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_956_inst flow-through 
    process(type_cast_956_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_956_inst:flowthrough inputs: " & " SUB_u2_u2_955_wire = "& Convert_SLV_To_Hex_String(SUB_u2_u2_955_wire) & " outputs:" & " type_cast_956_wire= "  & Convert_SLV_To_Hex_String(type_cast_956_wire));
      --
    end process; 
    -- interlock type_cast_956_inst
    process(SUB_u2_u2_955_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := SUB_u2_u2_955_wire(1 downto 0);
      type_cast_956_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_966_inst flow-through 
    process(type_cast_966_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_966_inst:flowthrough inputs: " & " SUB_u2_u2_965_wire = "& Convert_SLV_To_Hex_String(SUB_u2_u2_965_wire) & " outputs:" & " type_cast_966_wire= "  & Convert_SLV_To_Hex_String(type_cast_966_wire));
      --
    end process; 
    -- interlock type_cast_966_inst
    process(SUB_u2_u2_965_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := SUB_u2_u2_965_wire(1 downto 0);
      type_cast_966_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_970_inst flow-through 
    process(type_cast_970_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_970_inst:flowthrough inputs: " & " ADD_u2_u2_969_wire = "& Convert_SLV_To_Hex_String(ADD_u2_u2_969_wire) & " outputs:" & " type_cast_970_wire= "  & Convert_SLV_To_Hex_String(type_cast_970_wire));
      --
    end process; 
    -- interlock type_cast_970_inst
    process(ADD_u2_u2_969_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := ADD_u2_u2_969_wire(1 downto 0);
      type_cast_970_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_982_inst flow-through 
    process(type_cast_982_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_982_inst:flowthrough inputs: " & " ADD_u2_u2_981_wire = "& Convert_SLV_To_Hex_String(ADD_u2_u2_981_wire) & " outputs:" & " type_cast_982_wire= "  & Convert_SLV_To_Hex_String(type_cast_982_wire));
      --
    end process; 
    -- interlock type_cast_982_inst
    process(ADD_u2_u2_981_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := ADD_u2_u2_981_wire(1 downto 0);
      type_cast_982_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_993_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_993_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_993_inst:started:   inputs: " & " MUL_u16_u16_992_wire = "& Convert_SLV_To_Hex_String(MUL_u16_u16_992_wire));
          --
        end if; 
        if type_cast_993_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:type_cast_993_inst:finished:  outputs: " & " pp03_994= "  & Convert_SLV_To_Hex_String(pp03_994));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_993_inst_req_0;
      type_cast_993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_993_inst_req_1;
      type_cast_993_inst_ack_1<= rack(0);
      type_cast_993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        full_rate =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag => true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => MUL_u16_u16_992_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pp03_994,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_1001_gather_scatter flow-through 
    process(array_obj_ref_1001_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1001_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1001_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1001_data_0) & "outputs: " & " array_obj_ref_1001_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1001_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1001_gather_scatter
    process(array_obj_ref_1001_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1001_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1001_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1008_addr_0 flow-through 
    process(array_obj_ref_1008_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_addr_0:flowthrough  inputs: " & " array_obj_ref_1008_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_root_address) & "outputs: " & " array_obj_ref_1008_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1008_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1008_addr_0
    process(array_obj_ref_1008_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1008_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1008_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1008_gather_scatter flow-through 
    process(array_obj_ref_1008_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1008_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_data_0) & "outputs: " & " array_obj_ref_1008_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1008_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1008_gather_scatter
    process(array_obj_ref_1008_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1008_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1008_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1008_index_1_rename flow-through 
    process(R_col_to_be_replaced_1007_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1007_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1007_resized) & "outputs: " & " R_col_to_be_replaced_1007_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1007_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1008_index_1_rename
    process(R_col_to_be_replaced_1007_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1007_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1007_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1008_index_1_resize flow-through 
    process(R_col_to_be_replaced_1007_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_1007_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1007_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1008_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1007_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1008_root_address_inst flow-through 
    process(array_obj_ref_1008_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1008_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_final_offset) & "outputs: " & " array_obj_ref_1008_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1008_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1008_root_address_inst
    process(array_obj_ref_1008_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1008_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1008_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1011_gather_scatter flow-through 
    process(array_obj_ref_1011_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1011_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1011_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1011_data_0) & "outputs: " & " array_obj_ref_1011_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1011_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1011_gather_scatter
    process(array_obj_ref_1011_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1011_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1011_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1018_addr_0 flow-through 
    process(array_obj_ref_1018_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_addr_0:flowthrough  inputs: " & " array_obj_ref_1018_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_root_address) & "outputs: " & " array_obj_ref_1018_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1018_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1018_addr_0
    process(array_obj_ref_1018_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1018_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1018_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1018_gather_scatter flow-through 
    process(array_obj_ref_1018_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1018_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_data_0) & "outputs: " & " array_obj_ref_1018_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1018_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1018_gather_scatter
    process(array_obj_ref_1018_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1018_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1018_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1018_index_1_rename flow-through 
    process(R_col_to_be_replaced_1017_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1017_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1017_resized) & "outputs: " & " R_col_to_be_replaced_1017_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1017_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1018_index_1_rename
    process(R_col_to_be_replaced_1017_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1017_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1017_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1018_index_1_resize flow-through 
    process(R_col_to_be_replaced_1017_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_1017_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1017_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1018_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1017_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1018_root_address_inst flow-through 
    process(array_obj_ref_1018_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1018_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_final_offset) & "outputs: " & " array_obj_ref_1018_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1018_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1018_root_address_inst
    process(array_obj_ref_1018_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1018_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1018_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1021_gather_scatter flow-through 
    process(array_obj_ref_1021_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1021_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1021_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1021_data_0) & "outputs: " & " array_obj_ref_1021_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1021_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1021_gather_scatter
    process(array_obj_ref_1021_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1021_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1021_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1028_addr_0 flow-through 
    process(array_obj_ref_1028_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_addr_0:flowthrough  inputs: " & " array_obj_ref_1028_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_root_address) & "outputs: " & " array_obj_ref_1028_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1028_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1028_addr_0
    process(array_obj_ref_1028_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1028_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1028_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1028_gather_scatter flow-through 
    process(array_obj_ref_1028_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1028_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_data_0) & "outputs: " & " array_obj_ref_1028_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1028_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1028_gather_scatter
    process(array_obj_ref_1028_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1028_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1028_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1028_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_1027_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_1027_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1027_resized) & "outputs: " & " R_col_to_be_replaced_1_1027_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1027_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1028_index_1_rename
    process(R_col_to_be_replaced_1_1027_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_1027_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_1027_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1028_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_1027_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_958 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_958) & "outputs: " & " R_col_to_be_replaced_1_1027_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1027_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1028_index_1_resize
    process(col_to_be_replaced_1_958) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_958;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_1027_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1028_root_address_inst flow-through 
    process(array_obj_ref_1028_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1028_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_final_offset) & "outputs: " & " array_obj_ref_1028_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1028_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1028_root_address_inst
    process(array_obj_ref_1028_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1028_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1028_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1031_gather_scatter flow-through 
    process(array_obj_ref_1031_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1031_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1031_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1031_data_0) & "outputs: " & " array_obj_ref_1031_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1031_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1031_gather_scatter
    process(array_obj_ref_1031_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1031_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1031_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1038_addr_0 flow-through 
    process(array_obj_ref_1038_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_addr_0:flowthrough  inputs: " & " array_obj_ref_1038_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_root_address) & "outputs: " & " array_obj_ref_1038_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1038_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1038_addr_0
    process(array_obj_ref_1038_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1038_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1038_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1038_gather_scatter flow-through 
    process(array_obj_ref_1038_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1038_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_data_0) & "outputs: " & " array_obj_ref_1038_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1038_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1038_gather_scatter
    process(array_obj_ref_1038_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1038_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1038_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1038_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_1037_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_1037_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1037_resized) & "outputs: " & " R_col_to_be_replaced_1_1037_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1037_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1038_index_1_rename
    process(R_col_to_be_replaced_1_1037_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_1037_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_1037_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1038_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_1037_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_958 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_958) & "outputs: " & " R_col_to_be_replaced_1_1037_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1037_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1038_index_1_resize
    process(col_to_be_replaced_1_958) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_958;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_1037_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1038_root_address_inst flow-through 
    process(array_obj_ref_1038_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1038_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_final_offset) & "outputs: " & " array_obj_ref_1038_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1038_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1038_root_address_inst
    process(array_obj_ref_1038_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1038_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1038_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1041_gather_scatter flow-through 
    process(array_obj_ref_1041_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1041_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1041_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1041_data_0) & "outputs: " & " array_obj_ref_1041_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1041_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1041_gather_scatter
    process(array_obj_ref_1041_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1041_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1041_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1048_addr_0 flow-through 
    process(array_obj_ref_1048_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_addr_0:flowthrough  inputs: " & " array_obj_ref_1048_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_root_address) & "outputs: " & " array_obj_ref_1048_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1048_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1048_addr_0
    process(array_obj_ref_1048_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1048_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1048_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1048_gather_scatter flow-through 
    process(array_obj_ref_1048_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1048_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_data_0) & "outputs: " & " array_obj_ref_1048_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1048_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1048_gather_scatter
    process(array_obj_ref_1048_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1048_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1048_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1048_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_1047_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_1047_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1047_resized) & "outputs: " & " R_col_to_be_replaced_1_1047_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1047_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1048_index_1_rename
    process(R_col_to_be_replaced_1_1047_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_1047_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_1047_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1048_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_1047_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_958 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_958) & "outputs: " & " R_col_to_be_replaced_1_1047_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1047_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1048_index_1_resize
    process(col_to_be_replaced_1_958) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_958;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_1047_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1048_root_address_inst flow-through 
    process(array_obj_ref_1048_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1048_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_final_offset) & "outputs: " & " array_obj_ref_1048_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1048_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1048_root_address_inst
    process(array_obj_ref_1048_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1048_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1048_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1051_gather_scatter flow-through 
    process(array_obj_ref_1051_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1051_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1051_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1051_data_0) & "outputs: " & " array_obj_ref_1051_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1051_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1051_gather_scatter
    process(array_obj_ref_1051_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1051_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1051_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1058_addr_0 flow-through 
    process(array_obj_ref_1058_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_addr_0:flowthrough  inputs: " & " array_obj_ref_1058_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_root_address) & "outputs: " & " array_obj_ref_1058_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1058_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1058_addr_0
    process(array_obj_ref_1058_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1058_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1058_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1058_gather_scatter flow-through 
    process(array_obj_ref_1058_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1058_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_data_0) & "outputs: " & " array_obj_ref_1058_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1058_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1058_gather_scatter
    process(array_obj_ref_1058_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1058_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1058_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1058_index_1_rename flow-through 
    process(R_col_to_be_replaced_1_1057_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_1_1057_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1057_resized) & "outputs: " & " R_col_to_be_replaced_1_1057_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1057_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1058_index_1_rename
    process(R_col_to_be_replaced_1_1057_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_1_1057_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_1_1057_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1058_index_1_resize flow-through 
    process(R_col_to_be_replaced_1_1057_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_1_958 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_1_958) & "outputs: " & " R_col_to_be_replaced_1_1057_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1057_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1058_index_1_resize
    process(col_to_be_replaced_1_958) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_1_958;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_1_1057_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1058_root_address_inst flow-through 
    process(array_obj_ref_1058_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1058_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_final_offset) & "outputs: " & " array_obj_ref_1058_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1058_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1058_root_address_inst
    process(array_obj_ref_1058_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1058_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1058_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1061_gather_scatter flow-through 
    process(array_obj_ref_1061_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1061_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1061_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1061_data_0) & "outputs: " & " array_obj_ref_1061_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1061_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1061_gather_scatter
    process(array_obj_ref_1061_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1061_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1061_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1068_addr_0 flow-through 
    process(array_obj_ref_1068_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_addr_0:flowthrough  inputs: " & " array_obj_ref_1068_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_root_address) & "outputs: " & " array_obj_ref_1068_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1068_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1068_addr_0
    process(array_obj_ref_1068_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1068_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1068_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1068_gather_scatter flow-through 
    process(array_obj_ref_1068_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1068_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_data_0) & "outputs: " & " array_obj_ref_1068_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1068_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1068_gather_scatter
    process(array_obj_ref_1068_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1068_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1068_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1068_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_1067_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_1067_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1067_resized) & "outputs: " & " R_col_to_be_replaced_2_1067_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1067_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1068_index_1_rename
    process(R_col_to_be_replaced_2_1067_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_1067_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_1067_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1068_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_1067_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_972 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_972) & "outputs: " & " R_col_to_be_replaced_2_1067_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1067_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1068_index_1_resize
    process(col_to_be_replaced_2_972) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_972;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_1067_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1068_root_address_inst flow-through 
    process(array_obj_ref_1068_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1068_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_final_offset) & "outputs: " & " array_obj_ref_1068_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1068_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1068_root_address_inst
    process(array_obj_ref_1068_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1068_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1068_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1071_gather_scatter flow-through 
    process(array_obj_ref_1071_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1071_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1071_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1071_data_0) & "outputs: " & " array_obj_ref_1071_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1071_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1071_gather_scatter
    process(array_obj_ref_1071_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1071_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1071_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1078_addr_0 flow-through 
    process(array_obj_ref_1078_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_addr_0:flowthrough  inputs: " & " array_obj_ref_1078_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_root_address) & "outputs: " & " array_obj_ref_1078_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1078_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1078_addr_0
    process(array_obj_ref_1078_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1078_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1078_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1078_gather_scatter flow-through 
    process(array_obj_ref_1078_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1078_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_data_0) & "outputs: " & " array_obj_ref_1078_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1078_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1078_gather_scatter
    process(array_obj_ref_1078_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1078_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1078_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1078_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_1077_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_1077_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1077_resized) & "outputs: " & " R_col_to_be_replaced_2_1077_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1077_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1078_index_1_rename
    process(R_col_to_be_replaced_2_1077_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_1077_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_1077_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1078_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_1077_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_972 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_972) & "outputs: " & " R_col_to_be_replaced_2_1077_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1077_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1078_index_1_resize
    process(col_to_be_replaced_2_972) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_972;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_1077_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1078_root_address_inst flow-through 
    process(array_obj_ref_1078_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1078_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_final_offset) & "outputs: " & " array_obj_ref_1078_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1078_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1078_root_address_inst
    process(array_obj_ref_1078_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1078_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1078_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1081_gather_scatter flow-through 
    process(array_obj_ref_1081_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1081_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1081_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1081_data_0) & "outputs: " & " array_obj_ref_1081_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1081_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1081_gather_scatter
    process(array_obj_ref_1081_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1081_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1081_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1088_addr_0 flow-through 
    process(array_obj_ref_1088_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_addr_0:flowthrough  inputs: " & " array_obj_ref_1088_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_root_address) & "outputs: " & " array_obj_ref_1088_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1088_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1088_addr_0
    process(array_obj_ref_1088_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1088_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1088_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1088_gather_scatter flow-through 
    process(array_obj_ref_1088_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1088_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_data_0) & "outputs: " & " array_obj_ref_1088_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1088_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1088_gather_scatter
    process(array_obj_ref_1088_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1088_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1088_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1088_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_1087_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_1087_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1087_resized) & "outputs: " & " R_col_to_be_replaced_2_1087_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1087_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1088_index_1_rename
    process(R_col_to_be_replaced_2_1087_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_1087_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_1087_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1088_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_1087_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_972 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_972) & "outputs: " & " R_col_to_be_replaced_2_1087_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1087_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1088_index_1_resize
    process(col_to_be_replaced_2_972) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_972;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_1087_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1088_root_address_inst flow-through 
    process(array_obj_ref_1088_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1088_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_final_offset) & "outputs: " & " array_obj_ref_1088_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1088_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1088_root_address_inst
    process(array_obj_ref_1088_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1088_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1088_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1091_gather_scatter flow-through 
    process(array_obj_ref_1091_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1091_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1091_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1091_data_0) & "outputs: " & " array_obj_ref_1091_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1091_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1091_gather_scatter
    process(array_obj_ref_1091_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1091_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1091_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1098_addr_0 flow-through 
    process(array_obj_ref_1098_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_addr_0:flowthrough  inputs: " & " array_obj_ref_1098_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_root_address) & "outputs: " & " array_obj_ref_1098_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1098_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1098_addr_0
    process(array_obj_ref_1098_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1098_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1098_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1098_gather_scatter flow-through 
    process(array_obj_ref_1098_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1098_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_data_0) & "outputs: " & " array_obj_ref_1098_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1098_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1098_gather_scatter
    process(array_obj_ref_1098_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1098_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1098_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1098_index_1_rename flow-through 
    process(R_col_to_be_replaced_2_1097_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_2_1097_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1097_resized) & "outputs: " & " R_col_to_be_replaced_2_1097_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1097_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1098_index_1_rename
    process(R_col_to_be_replaced_2_1097_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_2_1097_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_2_1097_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1098_index_1_resize flow-through 
    process(R_col_to_be_replaced_2_1097_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_2_972 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_2_972) & "outputs: " & " R_col_to_be_replaced_2_1097_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1097_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1098_index_1_resize
    process(col_to_be_replaced_2_972) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_2_972;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_2_1097_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1098_root_address_inst flow-through 
    process(array_obj_ref_1098_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1098_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_final_offset) & "outputs: " & " array_obj_ref_1098_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1098_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1098_root_address_inst
    process(array_obj_ref_1098_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1098_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1098_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1101_gather_scatter flow-through 
    process(array_obj_ref_1101_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1101_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1101_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1101_data_0) & "outputs: " & " array_obj_ref_1101_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1101_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1101_gather_scatter
    process(array_obj_ref_1101_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1101_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1101_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1108_addr_0 flow-through 
    process(array_obj_ref_1108_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_addr_0:flowthrough  inputs: " & " array_obj_ref_1108_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_root_address) & "outputs: " & " array_obj_ref_1108_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1108_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1108_addr_0
    process(array_obj_ref_1108_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1108_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1108_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1108_gather_scatter flow-through 
    process(array_obj_ref_1108_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1108_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_data_0) & "outputs: " & " array_obj_ref_1108_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1108_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1108_gather_scatter
    process(array_obj_ref_1108_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1108_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1108_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1108_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_1107_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_1107_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1107_resized) & "outputs: " & " R_col_to_be_replaced_3_1107_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1107_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1108_index_1_rename
    process(R_col_to_be_replaced_3_1107_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_1107_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_1107_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1108_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_1107_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_984 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_984) & "outputs: " & " R_col_to_be_replaced_3_1107_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1107_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1108_index_1_resize
    process(col_to_be_replaced_3_984) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_984;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_1107_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1108_root_address_inst flow-through 
    process(array_obj_ref_1108_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1108_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_final_offset) & "outputs: " & " array_obj_ref_1108_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1108_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1108_root_address_inst
    process(array_obj_ref_1108_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1108_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1108_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1111_gather_scatter flow-through 
    process(array_obj_ref_1111_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1111_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1111_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1111_data_0) & "outputs: " & " array_obj_ref_1111_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1111_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1111_gather_scatter
    process(array_obj_ref_1111_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1111_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1111_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1118_addr_0 flow-through 
    process(array_obj_ref_1118_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_addr_0:flowthrough  inputs: " & " array_obj_ref_1118_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_root_address) & "outputs: " & " array_obj_ref_1118_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1118_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1118_addr_0
    process(array_obj_ref_1118_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1118_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1118_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1118_gather_scatter flow-through 
    process(array_obj_ref_1118_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1118_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_data_0) & "outputs: " & " array_obj_ref_1118_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1118_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1118_gather_scatter
    process(array_obj_ref_1118_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1118_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1118_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1118_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_1117_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_1117_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1117_resized) & "outputs: " & " R_col_to_be_replaced_3_1117_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1117_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1118_index_1_rename
    process(R_col_to_be_replaced_3_1117_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_1117_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_1117_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1118_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_1117_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_984 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_984) & "outputs: " & " R_col_to_be_replaced_3_1117_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1117_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1118_index_1_resize
    process(col_to_be_replaced_3_984) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_984;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_1117_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1118_root_address_inst flow-through 
    process(array_obj_ref_1118_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1118_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_final_offset) & "outputs: " & " array_obj_ref_1118_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1118_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1118_root_address_inst
    process(array_obj_ref_1118_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1118_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1118_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1121_gather_scatter flow-through 
    process(array_obj_ref_1121_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1121_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1121_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1121_data_0) & "outputs: " & " array_obj_ref_1121_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1121_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1121_gather_scatter
    process(array_obj_ref_1121_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1121_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1121_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1128_addr_0 flow-through 
    process(array_obj_ref_1128_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_addr_0:flowthrough  inputs: " & " array_obj_ref_1128_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_root_address) & "outputs: " & " array_obj_ref_1128_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1128_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1128_addr_0
    process(array_obj_ref_1128_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1128_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1128_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1128_gather_scatter flow-through 
    process(array_obj_ref_1128_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1128_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_data_0) & "outputs: " & " array_obj_ref_1128_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1128_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1128_gather_scatter
    process(array_obj_ref_1128_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1128_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1128_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1128_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_1127_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_1127_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1127_resized) & "outputs: " & " R_col_to_be_replaced_3_1127_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1127_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1128_index_1_rename
    process(R_col_to_be_replaced_3_1127_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_1127_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_1127_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1128_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_1127_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_984 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_984) & "outputs: " & " R_col_to_be_replaced_3_1127_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1127_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1128_index_1_resize
    process(col_to_be_replaced_3_984) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_984;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_1127_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1128_root_address_inst flow-through 
    process(array_obj_ref_1128_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1128_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_final_offset) & "outputs: " & " array_obj_ref_1128_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1128_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1128_root_address_inst
    process(array_obj_ref_1128_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1128_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1128_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1131_gather_scatter flow-through 
    process(array_obj_ref_1131_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1131_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1131_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1131_data_0) & "outputs: " & " array_obj_ref_1131_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1131_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1131_gather_scatter
    process(array_obj_ref_1131_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1131_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1131_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1138_addr_0 flow-through 
    process(array_obj_ref_1138_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_addr_0:flowthrough  inputs: " & " array_obj_ref_1138_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_root_address) & "outputs: " & " array_obj_ref_1138_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1138_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1138_addr_0
    process(array_obj_ref_1138_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1138_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_1138_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1138_gather_scatter flow-through 
    process(array_obj_ref_1138_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1138_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_data_0) & "outputs: " & " array_obj_ref_1138_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1138_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1138_gather_scatter
    process(array_obj_ref_1138_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1138_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1138_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1138_index_1_rename flow-through 
    process(R_col_to_be_replaced_3_1137_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_3_1137_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1137_resized) & "outputs: " & " R_col_to_be_replaced_3_1137_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1137_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1138_index_1_rename
    process(R_col_to_be_replaced_3_1137_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_3_1137_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_3_1137_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1138_index_1_resize flow-through 
    process(R_col_to_be_replaced_3_1137_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_3_984 = "& Convert_SLV_To_Hex_String(col_to_be_replaced_3_984) & "outputs: " & " R_col_to_be_replaced_3_1137_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1137_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1138_index_1_resize
    process(col_to_be_replaced_3_984) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_3_984;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_3_1137_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1138_root_address_inst flow-through 
    process(array_obj_ref_1138_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1138_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_final_offset) & "outputs: " & " array_obj_ref_1138_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1138_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1138_root_address_inst
    process(array_obj_ref_1138_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1138_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_1138_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1141_gather_scatter flow-through 
    process(array_obj_ref_1141_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1141_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1141_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1141_data_0) & "outputs: " & " array_obj_ref_1141_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1141_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1141_gather_scatter
    process(array_obj_ref_1141_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1141_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_1141_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_988_addr_0 flow-through 
    process(array_obj_ref_988_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_addr_0:flowthrough  inputs: " & " array_obj_ref_988_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_988_root_address) & "outputs: " & " array_obj_ref_988_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_988_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_988_addr_0
    process(array_obj_ref_988_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_988_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_988_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_988_gather_scatter flow-through 
    process(array_obj_ref_988_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_gather_scatter:flowthrough  inputs: " & " array_obj_ref_988_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_988_data_0) & "outputs: " & " array_obj_ref_988_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_988_wire));
      --
    end process; 
    -- equivalence array_obj_ref_988_gather_scatter
    process(array_obj_ref_988_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_988_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_988_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_988_index_1_rename flow-through 
    process(R_col_to_be_replaced_987_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_987_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_987_resized) & "outputs: " & " R_col_to_be_replaced_987_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_987_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_988_index_1_rename
    process(R_col_to_be_replaced_987_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_987_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_987_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_988_index_1_resize flow-through 
    process(R_col_to_be_replaced_987_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_987_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_987_resized));
      --
    end process; 
    -- equivalence array_obj_ref_988_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_987_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_988_root_address_inst flow-through 
    process(array_obj_ref_988_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_root_address_inst:flowthrough  inputs: " & " array_obj_ref_988_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_988_final_offset) & "outputs: " & " array_obj_ref_988_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_988_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_988_root_address_inst
    process(array_obj_ref_988_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_988_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_988_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_991_gather_scatter flow-through 
    process(array_obj_ref_991_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_991_gather_scatter:flowthrough  inputs: " & " array_obj_ref_991_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_991_data_0) & "outputs: " & " array_obj_ref_991_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_991_wire));
      --
    end process; 
    -- equivalence array_obj_ref_991_gather_scatter
    process(array_obj_ref_991_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_991_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_991_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_998_addr_0 flow-through 
    process(array_obj_ref_998_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_addr_0:flowthrough  inputs: " & " array_obj_ref_998_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_998_root_address) & "outputs: " & " array_obj_ref_998_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_998_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_998_addr_0
    process(array_obj_ref_998_root_address) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_998_root_address;
      ov(3 downto 0) := iv;
      array_obj_ref_998_word_address_0 <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_998_gather_scatter flow-through 
    process(array_obj_ref_998_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_gather_scatter:flowthrough  inputs: " & " array_obj_ref_998_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_998_data_0) & "outputs: " & " array_obj_ref_998_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_998_wire));
      --
    end process; 
    -- equivalence array_obj_ref_998_gather_scatter
    process(array_obj_ref_998_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_998_data_0;
      ov(15 downto 0) := iv;
      array_obj_ref_998_wire <= ov(15 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_998_index_1_rename flow-through 
    process(R_col_to_be_replaced_997_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_index_1_rename:flowthrough  inputs: " & " R_col_to_be_replaced_997_resized = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_997_resized) & "outputs: " & " R_col_to_be_replaced_997_scaled= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_997_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_998_index_1_rename
    process(R_col_to_be_replaced_997_resized) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_col_to_be_replaced_997_resized;
      ov(3 downto 0) := iv;
      R_col_to_be_replaced_997_scaled <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_998_index_1_resize flow-through 
    process(R_col_to_be_replaced_997_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_index_1_resize:flowthrough  inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & "outputs: " & " R_col_to_be_replaced_997_resized= "  & Convert_SLV_To_Hex_String(R_col_to_be_replaced_997_resized));
      --
    end process; 
    -- equivalence array_obj_ref_998_index_1_resize
    process(col_to_be_replaced_buffer) --
      variable iv : std_logic_vector(1 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := col_to_be_replaced_buffer;
      ov(1 downto 0) := iv;
      R_col_to_be_replaced_997_resized <= ov(3 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_998_root_address_inst flow-through 
    process(array_obj_ref_998_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_root_address_inst:flowthrough  inputs: " & " array_obj_ref_998_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_998_final_offset) & "outputs: " & " array_obj_ref_998_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_998_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_998_root_address_inst
    process(array_obj_ref_998_final_offset) --
      variable iv : std_logic_vector(3 downto 0);
      variable ov : std_logic_vector(3 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_998_final_offset;
      ov(3 downto 0) := iv;
      array_obj_ref_998_root_address <= ov(3 downto 0);
      --
    end process;
    -- logger for split-operator ADD_u16_u16_1148_inst flow-through 
    process(ADD_u16_u16_1148_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1148_inst:flowthrough inputs: " & " pp00_1114 = "& Convert_SLV_To_Hex_String(pp00_1114) & " pp01_1074 = "& Convert_SLV_To_Hex_String(pp01_1074) & " outputs:" & " ADD_u16_u16_1148_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1148_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1148_inst
    process(pp00_1114, pp01_1074) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp00_1114, pp01_1074, tmp_var);
      ADD_u16_u16_1148_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1154_inst flow-through 
    process(ADD_u16_u16_1154_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1154_inst:flowthrough inputs: " & " pp02_1034 = "& Convert_SLV_To_Hex_String(pp02_1034) & " pp03_994 = "& Convert_SLV_To_Hex_String(pp03_994) & " outputs:" & " ADD_u16_u16_1154_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1154_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1154_inst
    process(pp02_1034, pp03_994) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp02_1034, pp03_994, tmp_var);
      ADD_u16_u16_1154_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1160_inst flow-through 
    process(ADD_u16_u16_1160_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1160_inst:flowthrough inputs: " & " pp10_1124 = "& Convert_SLV_To_Hex_String(pp10_1124) & " pp11_1084 = "& Convert_SLV_To_Hex_String(pp11_1084) & " outputs:" & " ADD_u16_u16_1160_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1160_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1160_inst
    process(pp10_1124, pp11_1084) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp10_1124, pp11_1084, tmp_var);
      ADD_u16_u16_1160_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1166_inst flow-through 
    process(ADD_u16_u16_1166_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1166_inst:flowthrough inputs: " & " pp12_1044 = "& Convert_SLV_To_Hex_String(pp12_1044) & " pp13_1004 = "& Convert_SLV_To_Hex_String(pp13_1004) & " outputs:" & " ADD_u16_u16_1166_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1166_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1166_inst
    process(pp12_1044, pp13_1004) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp12_1044, pp13_1004, tmp_var);
      ADD_u16_u16_1166_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1172_inst flow-through 
    process(ADD_u16_u16_1172_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1172_inst:flowthrough inputs: " & " pp20_1134 = "& Convert_SLV_To_Hex_String(pp20_1134) & " pp21_1094 = "& Convert_SLV_To_Hex_String(pp21_1094) & " outputs:" & " ADD_u16_u16_1172_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1172_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1172_inst
    process(pp20_1134, pp21_1094) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp20_1134, pp21_1094, tmp_var);
      ADD_u16_u16_1172_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1178_inst flow-through 
    process(ADD_u16_u16_1178_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1178_inst:flowthrough inputs: " & " pp22_1054 = "& Convert_SLV_To_Hex_String(pp22_1054) & " pp23_1014 = "& Convert_SLV_To_Hex_String(pp23_1014) & " outputs:" & " ADD_u16_u16_1178_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1178_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1178_inst
    process(pp22_1054, pp23_1014) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp22_1054, pp23_1014, tmp_var);
      ADD_u16_u16_1178_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1184_inst flow-through 
    process(ADD_u16_u16_1184_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1184_inst:flowthrough inputs: " & " pp30_1144 = "& Convert_SLV_To_Hex_String(pp30_1144) & " pp31_1104 = "& Convert_SLV_To_Hex_String(pp31_1104) & " outputs:" & " ADD_u16_u16_1184_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1184_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1184_inst
    process(pp30_1144, pp31_1104) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp30_1144, pp31_1104, tmp_var);
      ADD_u16_u16_1184_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1190_inst flow-through 
    process(ADD_u16_u16_1190_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1190_inst:flowthrough inputs: " & " pp32_1064 = "& Convert_SLV_To_Hex_String(pp32_1064) & " pp33_1024 = "& Convert_SLV_To_Hex_String(pp33_1024) & " outputs:" & " ADD_u16_u16_1190_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1190_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1190_inst
    process(pp32_1064, pp33_1024) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pp32_1064, pp33_1024, tmp_var);
      ADD_u16_u16_1190_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1196_inst flow-through 
    process(ADD_u16_u16_1196_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1196_inst:flowthrough inputs: " & " sum0_1150 = "& Convert_SLV_To_Hex_String(sum0_1150) & " sum1_1156 = "& Convert_SLV_To_Hex_String(sum1_1156) & " outputs:" & " ADD_u16_u16_1196_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1196_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1196_inst
    process(sum0_1150, sum1_1156) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum0_1150, sum1_1156, tmp_var);
      ADD_u16_u16_1196_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1202_inst flow-through 
    process(ADD_u16_u16_1202_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1202_inst:flowthrough inputs: " & " sum2_1162 = "& Convert_SLV_To_Hex_String(sum2_1162) & " sum3_1168 = "& Convert_SLV_To_Hex_String(sum3_1168) & " outputs:" & " ADD_u16_u16_1202_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1202_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1202_inst
    process(sum2_1162, sum3_1168) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum2_1162, sum3_1168, tmp_var);
      ADD_u16_u16_1202_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1208_inst flow-through 
    process(ADD_u16_u16_1208_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1208_inst:flowthrough inputs: " & " sum4_1174 = "& Convert_SLV_To_Hex_String(sum4_1174) & " sum5_1180 = "& Convert_SLV_To_Hex_String(sum5_1180) & " outputs:" & " ADD_u16_u16_1208_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1208_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1208_inst
    process(sum4_1174, sum5_1180) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum4_1174, sum5_1180, tmp_var);
      ADD_u16_u16_1208_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1214_inst flow-through 
    process(ADD_u16_u16_1214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1214_inst:flowthrough inputs: " & " sum6_1186 = "& Convert_SLV_To_Hex_String(sum6_1186) & " sum7_1192 = "& Convert_SLV_To_Hex_String(sum7_1192) & " outputs:" & " ADD_u16_u16_1214_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1214_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1214_inst
    process(sum6_1186, sum7_1192) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum6_1186, sum7_1192, tmp_var);
      ADD_u16_u16_1214_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1220_inst flow-through 
    process(ADD_u16_u16_1220_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1220_inst:flowthrough inputs: " & " sum10_1198 = "& Convert_SLV_To_Hex_String(sum10_1198) & " sum11_1204 = "& Convert_SLV_To_Hex_String(sum11_1204) & " outputs:" & " ADD_u16_u16_1220_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1220_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1220_inst
    process(sum10_1198, sum11_1204) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum10_1198, sum11_1204, tmp_var);
      ADD_u16_u16_1220_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1226_inst flow-through 
    process(ADD_u16_u16_1226_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1226_inst:flowthrough inputs: " & " sum12_1210 = "& Convert_SLV_To_Hex_String(sum12_1210) & " sum13_1216 = "& Convert_SLV_To_Hex_String(sum13_1216) & " outputs:" & " ADD_u16_u16_1226_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1226_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1226_inst
    process(sum12_1210, sum13_1216) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum12_1210, sum13_1216, tmp_var);
      ADD_u16_u16_1226_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u16_u16_1232_inst flow-through 
    process(ADD_u16_u16_1232_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u16_u16_1232_inst:flowthrough inputs: " & " sum20_1222 = "& Convert_SLV_To_Hex_String(sum20_1222) & " sum21_1228 = "& Convert_SLV_To_Hex_String(sum21_1228) & " outputs:" & " ADD_u16_u16_1232_wire= "  & Convert_SLV_To_Hex_String(ADD_u16_u16_1232_wire));
      --
    end process; 
    -- binary operator ADD_u16_u16_1232_inst
    process(sum20_1222, sum21_1228) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sum20_1222, sum21_1228, tmp_var);
      ADD_u16_u16_1232_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u2_u2_969_inst flow-through 
    process(ADD_u2_u2_969_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u2_u2_969_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_968_wire_constant = "& Convert_SLV_To_Hex_String(konst_968_wire_constant) & " outputs:" & " ADD_u2_u2_969_wire= "  & Convert_SLV_To_Hex_String(ADD_u2_u2_969_wire));
      --
    end process; 
    -- binary operator ADD_u2_u2_969_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_to_be_replaced_buffer, konst_968_wire_constant, tmp_var);
      ADD_u2_u2_969_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u2_u2_981_inst flow-through 
    process(ADD_u2_u2_981_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:ADD_u2_u2_981_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_980_wire_constant = "& Convert_SLV_To_Hex_String(konst_980_wire_constant) & " outputs:" & " ADD_u2_u2_981_wire= "  & Convert_SLV_To_Hex_String(ADD_u2_u2_981_wire));
      --
    end process; 
    -- binary operator ADD_u2_u2_981_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_to_be_replaced_buffer, konst_980_wire_constant, tmp_var);
      ADD_u2_u2_981_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_950_inst flow-through 
    process(EQ_u2_u1_950_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:EQ_u2_u1_950_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_949_wire_constant = "& Convert_SLV_To_Hex_String(konst_949_wire_constant) & " outputs:" & " EQ_u2_u1_950_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_950_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_950_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_to_be_replaced_buffer, konst_949_wire_constant, tmp_var);
      EQ_u2_u1_950_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_976_inst flow-through 
    process(EQ_u2_u1_976_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:EQ_u2_u1_976_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_975_wire_constant = "& Convert_SLV_To_Hex_String(konst_975_wire_constant) & " outputs:" & " EQ_u2_u1_976_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_976_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_976_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_to_be_replaced_buffer, konst_975_wire_constant, tmp_var);
      EQ_u2_u1_976_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1002_inst flow-through 
    process(MUL_u16_u16_1002_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1002_inst:flowthrough inputs: " & " array_obj_ref_998_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_998_wire) & " array_obj_ref_1001_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1001_wire) & " outputs:" & " MUL_u16_u16_1002_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1002_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1002_inst
    process(array_obj_ref_998_wire, array_obj_ref_1001_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_998_wire, array_obj_ref_1001_wire, tmp_var);
      MUL_u16_u16_1002_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1012_inst flow-through 
    process(MUL_u16_u16_1012_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1012_inst:flowthrough inputs: " & " array_obj_ref_1008_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_wire) & " array_obj_ref_1011_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1011_wire) & " outputs:" & " MUL_u16_u16_1012_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1012_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1012_inst
    process(array_obj_ref_1008_wire, array_obj_ref_1011_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1008_wire, array_obj_ref_1011_wire, tmp_var);
      MUL_u16_u16_1012_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1022_inst flow-through 
    process(MUL_u16_u16_1022_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1022_inst:flowthrough inputs: " & " array_obj_ref_1018_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_wire) & " array_obj_ref_1021_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1021_wire) & " outputs:" & " MUL_u16_u16_1022_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1022_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1022_inst
    process(array_obj_ref_1018_wire, array_obj_ref_1021_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1018_wire, array_obj_ref_1021_wire, tmp_var);
      MUL_u16_u16_1022_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1032_inst flow-through 
    process(MUL_u16_u16_1032_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1032_inst:flowthrough inputs: " & " array_obj_ref_1028_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_wire) & " array_obj_ref_1031_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1031_wire) & " outputs:" & " MUL_u16_u16_1032_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1032_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1032_inst
    process(array_obj_ref_1028_wire, array_obj_ref_1031_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1028_wire, array_obj_ref_1031_wire, tmp_var);
      MUL_u16_u16_1032_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1042_inst flow-through 
    process(MUL_u16_u16_1042_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1042_inst:flowthrough inputs: " & " array_obj_ref_1038_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_wire) & " array_obj_ref_1041_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1041_wire) & " outputs:" & " MUL_u16_u16_1042_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1042_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1042_inst
    process(array_obj_ref_1038_wire, array_obj_ref_1041_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1038_wire, array_obj_ref_1041_wire, tmp_var);
      MUL_u16_u16_1042_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1052_inst flow-through 
    process(MUL_u16_u16_1052_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1052_inst:flowthrough inputs: " & " array_obj_ref_1048_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_wire) & " array_obj_ref_1051_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1051_wire) & " outputs:" & " MUL_u16_u16_1052_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1052_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1052_inst
    process(array_obj_ref_1048_wire, array_obj_ref_1051_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1048_wire, array_obj_ref_1051_wire, tmp_var);
      MUL_u16_u16_1052_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1062_inst flow-through 
    process(MUL_u16_u16_1062_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1062_inst:flowthrough inputs: " & " array_obj_ref_1058_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_wire) & " array_obj_ref_1061_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1061_wire) & " outputs:" & " MUL_u16_u16_1062_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1062_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1062_inst
    process(array_obj_ref_1058_wire, array_obj_ref_1061_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1058_wire, array_obj_ref_1061_wire, tmp_var);
      MUL_u16_u16_1062_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1072_inst flow-through 
    process(MUL_u16_u16_1072_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1072_inst:flowthrough inputs: " & " array_obj_ref_1068_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_wire) & " array_obj_ref_1071_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1071_wire) & " outputs:" & " MUL_u16_u16_1072_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1072_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1072_inst
    process(array_obj_ref_1068_wire, array_obj_ref_1071_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1068_wire, array_obj_ref_1071_wire, tmp_var);
      MUL_u16_u16_1072_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1082_inst flow-through 
    process(MUL_u16_u16_1082_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1082_inst:flowthrough inputs: " & " array_obj_ref_1078_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_wire) & " array_obj_ref_1081_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1081_wire) & " outputs:" & " MUL_u16_u16_1082_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1082_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1082_inst
    process(array_obj_ref_1078_wire, array_obj_ref_1081_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1078_wire, array_obj_ref_1081_wire, tmp_var);
      MUL_u16_u16_1082_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1092_inst flow-through 
    process(MUL_u16_u16_1092_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1092_inst:flowthrough inputs: " & " array_obj_ref_1088_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_wire) & " array_obj_ref_1091_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1091_wire) & " outputs:" & " MUL_u16_u16_1092_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1092_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1092_inst
    process(array_obj_ref_1088_wire, array_obj_ref_1091_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1088_wire, array_obj_ref_1091_wire, tmp_var);
      MUL_u16_u16_1092_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1102_inst flow-through 
    process(MUL_u16_u16_1102_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1102_inst:flowthrough inputs: " & " array_obj_ref_1098_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_wire) & " array_obj_ref_1101_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1101_wire) & " outputs:" & " MUL_u16_u16_1102_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1102_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1102_inst
    process(array_obj_ref_1098_wire, array_obj_ref_1101_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1098_wire, array_obj_ref_1101_wire, tmp_var);
      MUL_u16_u16_1102_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1112_inst flow-through 
    process(MUL_u16_u16_1112_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1112_inst:flowthrough inputs: " & " array_obj_ref_1108_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_wire) & " array_obj_ref_1111_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1111_wire) & " outputs:" & " MUL_u16_u16_1112_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1112_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1112_inst
    process(array_obj_ref_1108_wire, array_obj_ref_1111_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1108_wire, array_obj_ref_1111_wire, tmp_var);
      MUL_u16_u16_1112_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1122_inst flow-through 
    process(MUL_u16_u16_1122_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1122_inst:flowthrough inputs: " & " array_obj_ref_1118_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_wire) & " array_obj_ref_1121_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1121_wire) & " outputs:" & " MUL_u16_u16_1122_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1122_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1122_inst
    process(array_obj_ref_1118_wire, array_obj_ref_1121_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1118_wire, array_obj_ref_1121_wire, tmp_var);
      MUL_u16_u16_1122_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1132_inst flow-through 
    process(MUL_u16_u16_1132_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1132_inst:flowthrough inputs: " & " array_obj_ref_1128_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_wire) & " array_obj_ref_1131_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1131_wire) & " outputs:" & " MUL_u16_u16_1132_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1132_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1132_inst
    process(array_obj_ref_1128_wire, array_obj_ref_1131_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1128_wire, array_obj_ref_1131_wire, tmp_var);
      MUL_u16_u16_1132_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_1142_inst flow-through 
    process(MUL_u16_u16_1142_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_1142_inst:flowthrough inputs: " & " array_obj_ref_1138_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_wire) & " array_obj_ref_1141_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1141_wire) & " outputs:" & " MUL_u16_u16_1142_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_1142_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_1142_inst
    process(array_obj_ref_1138_wire, array_obj_ref_1141_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_1138_wire, array_obj_ref_1141_wire, tmp_var);
      MUL_u16_u16_1142_wire <= tmp_var; --
    end process;
    -- logger for split-operator MUL_u16_u16_992_inst flow-through 
    process(MUL_u16_u16_992_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:MUL_u16_u16_992_inst:flowthrough inputs: " & " array_obj_ref_988_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_988_wire) & " array_obj_ref_991_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_991_wire) & " outputs:" & " MUL_u16_u16_992_wire= "  & Convert_SLV_To_Hex_String(MUL_u16_u16_992_wire));
      --
    end process; 
    -- binary operator MUL_u16_u16_992_inst
    process(array_obj_ref_988_wire, array_obj_ref_991_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(array_obj_ref_988_wire, array_obj_ref_991_wire, tmp_var);
      MUL_u16_u16_992_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u2_u2_955_inst flow-through 
    process(SUB_u2_u2_955_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:SUB_u2_u2_955_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_954_wire_constant = "& Convert_SLV_To_Hex_String(konst_954_wire_constant) & " outputs:" & " SUB_u2_u2_955_wire= "  & Convert_SLV_To_Hex_String(SUB_u2_u2_955_wire));
      --
    end process; 
    -- binary operator SUB_u2_u2_955_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntSub_proc(col_to_be_replaced_buffer, konst_954_wire_constant, tmp_var);
      SUB_u2_u2_955_wire <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u2_u2_965_inst flow-through 
    process(SUB_u2_u2_965_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:SUB_u2_u2_965_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_964_wire_constant = "& Convert_SLV_To_Hex_String(konst_964_wire_constant) & " outputs:" & " SUB_u2_u2_965_wire= "  & Convert_SLV_To_Hex_String(SUB_u2_u2_965_wire));
      --
    end process; 
    -- binary operator SUB_u2_u2_965_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntSub_proc(col_to_be_replaced_buffer, konst_964_wire_constant, tmp_var);
      SUB_u2_u2_965_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGE_u2_u1_962_inst flow-through 
    process(UGE_u2_u1_962_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:UGE_u2_u1_962_inst:flowthrough inputs: " & " col_to_be_replaced_buffer = "& Convert_SLV_To_Hex_String(col_to_be_replaced_buffer) & " konst_961_wire_constant = "& Convert_SLV_To_Hex_String(konst_961_wire_constant) & " outputs:" & " UGE_u2_u1_962_wire= "  & Convert_SLV_To_Hex_String(UGE_u2_u1_962_wire));
      --
    end process; 
    -- binary operator UGE_u2_u1_962_inst
    process(col_to_be_replaced_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(col_to_be_replaced_buffer, konst_961_wire_constant, tmp_var);
      UGE_u2_u1_962_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_1008_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1008_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_index_offset:started:   inputs: " & " R_col_to_be_replaced_1007_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1007_scaled) & " array_obj_ref_1008_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1008_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_index_offset:finished:  outputs: " & " array_obj_ref_1008_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1008_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (38) : array_obj_ref_1008_index_offset 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1007_scaled;
      array_obj_ref_1008_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1008_index_offset_req_0;
      array_obj_ref_1008_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1008_index_offset_req_1;
      array_obj_ref_1008_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- logger for split-operator array_obj_ref_1018_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1018_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_index_offset:started:   inputs: " & " R_col_to_be_replaced_1017_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1017_scaled) & " array_obj_ref_1018_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1018_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_index_offset:finished:  outputs: " & " array_obj_ref_1018_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1018_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (39) : array_obj_ref_1018_index_offset 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1017_scaled;
      array_obj_ref_1018_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1018_index_offset_req_0;
      array_obj_ref_1018_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1018_index_offset_req_1;
      array_obj_ref_1018_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_39_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- logger for split-operator array_obj_ref_1028_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1028_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_1027_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1027_scaled) & " array_obj_ref_1028_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1028_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_index_offset:finished:  outputs: " & " array_obj_ref_1028_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1028_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (40) : array_obj_ref_1028_index_offset 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_1027_scaled;
      array_obj_ref_1028_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1028_index_offset_req_0;
      array_obj_ref_1028_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1028_index_offset_req_1;
      array_obj_ref_1028_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_40_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_40_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_40",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- logger for split-operator array_obj_ref_1038_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1038_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_1037_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1037_scaled) & " array_obj_ref_1038_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1038_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_index_offset:finished:  outputs: " & " array_obj_ref_1038_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1038_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (41) : array_obj_ref_1038_index_offset 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_1037_scaled;
      array_obj_ref_1038_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1038_index_offset_req_0;
      array_obj_ref_1038_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1038_index_offset_req_1;
      array_obj_ref_1038_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- logger for split-operator array_obj_ref_1048_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1048_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_1047_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1047_scaled) & " array_obj_ref_1048_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1048_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_index_offset:finished:  outputs: " & " array_obj_ref_1048_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1048_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (42) : array_obj_ref_1048_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_1047_scaled;
      array_obj_ref_1048_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1048_index_offset_req_0;
      array_obj_ref_1048_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1048_index_offset_req_1;
      array_obj_ref_1048_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- logger for split-operator array_obj_ref_1058_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1058_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_index_offset:started:   inputs: " & " R_col_to_be_replaced_1_1057_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_1_1057_scaled) & " array_obj_ref_1058_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1058_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_index_offset:finished:  outputs: " & " array_obj_ref_1058_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1058_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (43) : array_obj_ref_1058_index_offset 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_1_1057_scaled;
      array_obj_ref_1058_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1058_index_offset_req_0;
      array_obj_ref_1058_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1058_index_offset_req_1;
      array_obj_ref_1058_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- logger for split-operator array_obj_ref_1068_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1068_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_1067_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1067_scaled) & " array_obj_ref_1068_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1068_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_index_offset:finished:  outputs: " & " array_obj_ref_1068_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1068_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (44) : array_obj_ref_1068_index_offset 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_1067_scaled;
      array_obj_ref_1068_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1068_index_offset_req_0;
      array_obj_ref_1068_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1068_index_offset_req_1;
      array_obj_ref_1068_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- logger for split-operator array_obj_ref_1078_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1078_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_1077_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1077_scaled) & " array_obj_ref_1078_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1078_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_index_offset:finished:  outputs: " & " array_obj_ref_1078_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1078_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (45) : array_obj_ref_1078_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_1077_scaled;
      array_obj_ref_1078_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1078_index_offset_req_0;
      array_obj_ref_1078_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1078_index_offset_req_1;
      array_obj_ref_1078_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- logger for split-operator array_obj_ref_1088_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1088_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_1087_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1087_scaled) & " array_obj_ref_1088_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1088_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_index_offset:finished:  outputs: " & " array_obj_ref_1088_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1088_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (46) : array_obj_ref_1088_index_offset 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_1087_scaled;
      array_obj_ref_1088_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1088_index_offset_req_0;
      array_obj_ref_1088_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1088_index_offset_req_1;
      array_obj_ref_1088_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_46_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- logger for split-operator array_obj_ref_1098_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1098_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_index_offset:started:   inputs: " & " R_col_to_be_replaced_2_1097_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_2_1097_scaled) & " array_obj_ref_1098_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1098_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_index_offset:finished:  outputs: " & " array_obj_ref_1098_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1098_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (47) : array_obj_ref_1098_index_offset 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_2_1097_scaled;
      array_obj_ref_1098_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1098_index_offset_req_0;
      array_obj_ref_1098_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1098_index_offset_req_1;
      array_obj_ref_1098_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_47_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_47_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_47",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- logger for split-operator array_obj_ref_1108_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1108_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_1107_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1107_scaled) & " array_obj_ref_1108_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1108_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_index_offset:finished:  outputs: " & " array_obj_ref_1108_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1108_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (48) : array_obj_ref_1108_index_offset 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_1107_scaled;
      array_obj_ref_1108_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1108_index_offset_req_0;
      array_obj_ref_1108_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1108_index_offset_req_1;
      array_obj_ref_1108_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_48_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_48_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_48",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- logger for split-operator array_obj_ref_1118_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1118_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_1117_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1117_scaled) & " array_obj_ref_1118_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1118_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_index_offset:finished:  outputs: " & " array_obj_ref_1118_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1118_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (49) : array_obj_ref_1118_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_1117_scaled;
      array_obj_ref_1118_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1118_index_offset_req_0;
      array_obj_ref_1118_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1118_index_offset_req_1;
      array_obj_ref_1118_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- logger for split-operator array_obj_ref_1128_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1128_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_1127_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1127_scaled) & " array_obj_ref_1128_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1128_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_index_offset:finished:  outputs: " & " array_obj_ref_1128_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1128_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (50) : array_obj_ref_1128_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_1127_scaled;
      array_obj_ref_1128_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1128_index_offset_req_0;
      array_obj_ref_1128_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1128_index_offset_req_1;
      array_obj_ref_1128_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- logger for split-operator array_obj_ref_1138_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1138_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_index_offset:started:   inputs: " & " R_col_to_be_replaced_3_1137_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_3_1137_scaled) & " array_obj_ref_1138_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_1138_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_index_offset:finished:  outputs: " & " array_obj_ref_1138_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1138_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (51) : array_obj_ref_1138_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_3_1137_scaled;
      array_obj_ref_1138_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1138_index_offset_req_0;
      array_obj_ref_1138_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1138_index_offset_req_1;
      array_obj_ref_1138_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "1100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- logger for split-operator array_obj_ref_988_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_988_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_index_offset:started:   inputs: " & " R_col_to_be_replaced_987_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_987_scaled) & " array_obj_ref_988_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_988_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_988_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_index_offset:finished:  outputs: " & " array_obj_ref_988_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_988_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (52) : array_obj_ref_988_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_987_scaled;
      array_obj_ref_988_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_988_index_offset_req_0;
      array_obj_ref_988_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_988_index_offset_req_1;
      array_obj_ref_988_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- logger for split-operator array_obj_ref_998_index_offset
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_998_index_offset_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_index_offset:started:   inputs: " & " R_col_to_be_replaced_997_scaled = "& Convert_SLV_To_Hex_String(R_col_to_be_replaced_997_scaled) & " array_obj_ref_998_constant_part_of_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_998_constant_part_of_offset));
          --
        end if; 
        if array_obj_ref_998_index_offset_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_index_offset:finished:  outputs: " & " array_obj_ref_998_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_998_final_offset));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (53) : array_obj_ref_998_index_offset 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_col_to_be_replaced_997_scaled;
      array_obj_ref_998_final_offset <= data_out(3 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_998_index_offset_req_0;
      array_obj_ref_998_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_998_index_offset_req_1;
      array_obj_ref_998_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0100",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- logger for split-operator array_obj_ref_1141_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1141_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1141_load_0:started:   inputs: " & " array_obj_ref_1141_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1141_word_address_0));
          --
        end if; 
        if array_obj_ref_1141_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1141_load_0:finished:  outputs: " & " array_obj_ref_1141_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1141_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_991_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_991_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_991_load_0:started:   inputs: " & " array_obj_ref_991_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_991_word_address_0));
          --
        end if; 
        if array_obj_ref_991_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_991_load_0:finished:  outputs: " & " array_obj_ref_991_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_991_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1011_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1011_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1011_load_0:started:   inputs: " & " array_obj_ref_1011_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1011_word_address_0));
          --
        end if; 
        if array_obj_ref_1011_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1011_load_0:finished:  outputs: " & " array_obj_ref_1011_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1011_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1001_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1001_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1001_load_0:started:   inputs: " & " array_obj_ref_1001_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1001_word_address_0));
          --
        end if; 
        if array_obj_ref_1001_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1001_load_0:finished:  outputs: " & " array_obj_ref_1001_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1001_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1021_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1021_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1021_load_0:started:   inputs: " & " array_obj_ref_1021_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1021_word_address_0));
          --
        end if; 
        if array_obj_ref_1021_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1021_load_0:finished:  outputs: " & " array_obj_ref_1021_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1021_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1031_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1031_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1031_load_0:started:   inputs: " & " array_obj_ref_1031_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1031_word_address_0));
          --
        end if; 
        if array_obj_ref_1031_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1031_load_0:finished:  outputs: " & " array_obj_ref_1031_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1031_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1041_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1041_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1041_load_0:started:   inputs: " & " array_obj_ref_1041_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1041_word_address_0));
          --
        end if; 
        if array_obj_ref_1041_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1041_load_0:finished:  outputs: " & " array_obj_ref_1041_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1041_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1051_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1051_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1051_load_0:started:   inputs: " & " array_obj_ref_1051_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1051_word_address_0));
          --
        end if; 
        if array_obj_ref_1051_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1051_load_0:finished:  outputs: " & " array_obj_ref_1051_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1051_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1061_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1061_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1061_load_0:started:   inputs: " & " array_obj_ref_1061_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1061_word_address_0));
          --
        end if; 
        if array_obj_ref_1061_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1061_load_0:finished:  outputs: " & " array_obj_ref_1061_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1061_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1071_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1071_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1071_load_0:started:   inputs: " & " array_obj_ref_1071_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1071_word_address_0));
          --
        end if; 
        if array_obj_ref_1071_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1071_load_0:finished:  outputs: " & " array_obj_ref_1071_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1071_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1081_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1081_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1081_load_0:started:   inputs: " & " array_obj_ref_1081_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1081_word_address_0));
          --
        end if; 
        if array_obj_ref_1081_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1081_load_0:finished:  outputs: " & " array_obj_ref_1081_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1081_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1091_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1091_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1091_load_0:started:   inputs: " & " array_obj_ref_1091_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1091_word_address_0));
          --
        end if; 
        if array_obj_ref_1091_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1091_load_0:finished:  outputs: " & " array_obj_ref_1091_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1091_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1101_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1101_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1101_load_0:started:   inputs: " & " array_obj_ref_1101_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1101_word_address_0));
          --
        end if; 
        if array_obj_ref_1101_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1101_load_0:finished:  outputs: " & " array_obj_ref_1101_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1101_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1111_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1111_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1111_load_0:started:   inputs: " & " array_obj_ref_1111_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1111_word_address_0));
          --
        end if; 
        if array_obj_ref_1111_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1111_load_0:finished:  outputs: " & " array_obj_ref_1111_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1111_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1121_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1121_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1121_load_0:started:   inputs: " & " array_obj_ref_1121_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1121_word_address_0));
          --
        end if; 
        if array_obj_ref_1121_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1121_load_0:finished:  outputs: " & " array_obj_ref_1121_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1121_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1131_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1131_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1131_load_0:started:   inputs: " & " array_obj_ref_1131_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1131_word_address_0));
          --
        end if; 
        if array_obj_ref_1131_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1131_load_0:finished:  outputs: " & " array_obj_ref_1131_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1131_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_1141_load_0 array_obj_ref_991_load_0 array_obj_ref_1011_load_0 array_obj_ref_1001_load_0 array_obj_ref_1021_load_0 array_obj_ref_1031_load_0 array_obj_ref_1041_load_0 array_obj_ref_1051_load_0 array_obj_ref_1061_load_0 array_obj_ref_1071_load_0 array_obj_ref_1081_load_0 array_obj_ref_1091_load_0 array_obj_ref_1101_load_0 array_obj_ref_1111_load_0 array_obj_ref_1121_load_0 array_obj_ref_1131_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1141_load_0_req_0,
        array_obj_ref_1141_load_0_ack_0,
        array_obj_ref_1141_load_0_req_1,
        array_obj_ref_1141_load_0_ack_1,
        "array_obj_ref_1141_load_0",
        "memory_space_0" ,
        array_obj_ref_1141_data_0,
        array_obj_ref_1141_word_address_0,
        "array_obj_ref_1141_data_0",
        "array_obj_ref_1141_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_991_load_0_req_0,
        array_obj_ref_991_load_0_ack_0,
        array_obj_ref_991_load_0_req_1,
        array_obj_ref_991_load_0_ack_1,
        "array_obj_ref_991_load_0",
        "memory_space_0" ,
        array_obj_ref_991_data_0,
        array_obj_ref_991_word_address_0,
        "array_obj_ref_991_data_0",
        "array_obj_ref_991_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1011_load_0_req_0,
        array_obj_ref_1011_load_0_ack_0,
        array_obj_ref_1011_load_0_req_1,
        array_obj_ref_1011_load_0_ack_1,
        "array_obj_ref_1011_load_0",
        "memory_space_0" ,
        array_obj_ref_1011_data_0,
        array_obj_ref_1011_word_address_0,
        "array_obj_ref_1011_data_0",
        "array_obj_ref_1011_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1001_load_0_req_0,
        array_obj_ref_1001_load_0_ack_0,
        array_obj_ref_1001_load_0_req_1,
        array_obj_ref_1001_load_0_ack_1,
        "array_obj_ref_1001_load_0",
        "memory_space_0" ,
        array_obj_ref_1001_data_0,
        array_obj_ref_1001_word_address_0,
        "array_obj_ref_1001_data_0",
        "array_obj_ref_1001_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1021_load_0_req_0,
        array_obj_ref_1021_load_0_ack_0,
        array_obj_ref_1021_load_0_req_1,
        array_obj_ref_1021_load_0_ack_1,
        "array_obj_ref_1021_load_0",
        "memory_space_0" ,
        array_obj_ref_1021_data_0,
        array_obj_ref_1021_word_address_0,
        "array_obj_ref_1021_data_0",
        "array_obj_ref_1021_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1031_load_0_req_0,
        array_obj_ref_1031_load_0_ack_0,
        array_obj_ref_1031_load_0_req_1,
        array_obj_ref_1031_load_0_ack_1,
        "array_obj_ref_1031_load_0",
        "memory_space_0" ,
        array_obj_ref_1031_data_0,
        array_obj_ref_1031_word_address_0,
        "array_obj_ref_1031_data_0",
        "array_obj_ref_1031_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1041_load_0_req_0,
        array_obj_ref_1041_load_0_ack_0,
        array_obj_ref_1041_load_0_req_1,
        array_obj_ref_1041_load_0_ack_1,
        "array_obj_ref_1041_load_0",
        "memory_space_0" ,
        array_obj_ref_1041_data_0,
        array_obj_ref_1041_word_address_0,
        "array_obj_ref_1041_data_0",
        "array_obj_ref_1041_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1051_load_0_req_0,
        array_obj_ref_1051_load_0_ack_0,
        array_obj_ref_1051_load_0_req_1,
        array_obj_ref_1051_load_0_ack_1,
        "array_obj_ref_1051_load_0",
        "memory_space_0" ,
        array_obj_ref_1051_data_0,
        array_obj_ref_1051_word_address_0,
        "array_obj_ref_1051_data_0",
        "array_obj_ref_1051_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1061_load_0_req_0,
        array_obj_ref_1061_load_0_ack_0,
        array_obj_ref_1061_load_0_req_1,
        array_obj_ref_1061_load_0_ack_1,
        "array_obj_ref_1061_load_0",
        "memory_space_0" ,
        array_obj_ref_1061_data_0,
        array_obj_ref_1061_word_address_0,
        "array_obj_ref_1061_data_0",
        "array_obj_ref_1061_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1071_load_0_req_0,
        array_obj_ref_1071_load_0_ack_0,
        array_obj_ref_1071_load_0_req_1,
        array_obj_ref_1071_load_0_ack_1,
        "array_obj_ref_1071_load_0",
        "memory_space_0" ,
        array_obj_ref_1071_data_0,
        array_obj_ref_1071_word_address_0,
        "array_obj_ref_1071_data_0",
        "array_obj_ref_1071_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1081_load_0_req_0,
        array_obj_ref_1081_load_0_ack_0,
        array_obj_ref_1081_load_0_req_1,
        array_obj_ref_1081_load_0_ack_1,
        "array_obj_ref_1081_load_0",
        "memory_space_0" ,
        array_obj_ref_1081_data_0,
        array_obj_ref_1081_word_address_0,
        "array_obj_ref_1081_data_0",
        "array_obj_ref_1081_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1091_load_0_req_0,
        array_obj_ref_1091_load_0_ack_0,
        array_obj_ref_1091_load_0_req_1,
        array_obj_ref_1091_load_0_ack_1,
        "array_obj_ref_1091_load_0",
        "memory_space_0" ,
        array_obj_ref_1091_data_0,
        array_obj_ref_1091_word_address_0,
        "array_obj_ref_1091_data_0",
        "array_obj_ref_1091_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1101_load_0_req_0,
        array_obj_ref_1101_load_0_ack_0,
        array_obj_ref_1101_load_0_req_1,
        array_obj_ref_1101_load_0_ack_1,
        "array_obj_ref_1101_load_0",
        "memory_space_0" ,
        array_obj_ref_1101_data_0,
        array_obj_ref_1101_word_address_0,
        "array_obj_ref_1101_data_0",
        "array_obj_ref_1101_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1111_load_0_req_0,
        array_obj_ref_1111_load_0_ack_0,
        array_obj_ref_1111_load_0_req_1,
        array_obj_ref_1111_load_0_ack_1,
        "array_obj_ref_1111_load_0",
        "memory_space_0" ,
        array_obj_ref_1111_data_0,
        array_obj_ref_1111_word_address_0,
        "array_obj_ref_1111_data_0",
        "array_obj_ref_1111_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1121_load_0_req_0,
        array_obj_ref_1121_load_0_ack_0,
        array_obj_ref_1121_load_0_req_1,
        array_obj_ref_1121_load_0_ack_1,
        "array_obj_ref_1121_load_0",
        "memory_space_0" ,
        array_obj_ref_1121_data_0,
        array_obj_ref_1121_word_address_0,
        "array_obj_ref_1121_data_0",
        "array_obj_ref_1121_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1131_load_0_req_0,
        array_obj_ref_1131_load_0_ack_0,
        array_obj_ref_1131_load_0_req_1,
        array_obj_ref_1131_load_0_ack_1,
        "array_obj_ref_1131_load_0",
        "memory_space_0" ,
        array_obj_ref_1131_data_0,
        array_obj_ref_1131_word_address_0,
        "array_obj_ref_1131_data_0",
        "array_obj_ref_1131_word_address_0" -- 
      );
      reqL_unguarded(15) <= array_obj_ref_1141_load_0_req_0;
      reqL_unguarded(14) <= array_obj_ref_991_load_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_1011_load_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_1001_load_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_1021_load_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_1031_load_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_1041_load_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_1051_load_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_1061_load_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_1071_load_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_1081_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_1091_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1101_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1111_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1121_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1131_load_0_req_0;
      array_obj_ref_1141_load_0_ack_0 <= ackL_unguarded(15);
      array_obj_ref_991_load_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_1011_load_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_1001_load_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_1021_load_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_1031_load_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_1041_load_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_1051_load_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_1061_load_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_1071_load_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_1081_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_1091_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1101_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1111_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1121_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1131_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= array_obj_ref_1141_load_0_req_1;
      reqR_unguarded(14) <= array_obj_ref_991_load_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_1011_load_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_1001_load_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_1021_load_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_1031_load_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_1041_load_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_1051_load_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_1061_load_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_1071_load_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_1081_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_1091_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1101_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1111_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1121_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1131_load_0_req_1;
      array_obj_ref_1141_load_0_ack_1 <= ackR_unguarded(15);
      array_obj_ref_991_load_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_1011_load_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_1001_load_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_1021_load_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_1031_load_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_1041_load_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_1051_load_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_1061_load_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_1071_load_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_1081_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_1091_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1101_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1111_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1121_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1131_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_15: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1141_word_address_0 & array_obj_ref_991_word_address_0 & array_obj_ref_1011_word_address_0 & array_obj_ref_1001_word_address_0 & array_obj_ref_1021_word_address_0 & array_obj_ref_1031_word_address_0 & array_obj_ref_1041_word_address_0 & array_obj_ref_1051_word_address_0 & array_obj_ref_1061_word_address_0 & array_obj_ref_1071_word_address_0 & array_obj_ref_1081_word_address_0 & array_obj_ref_1091_word_address_0 & array_obj_ref_1101_word_address_0 & array_obj_ref_1111_word_address_0 & array_obj_ref_1121_word_address_0 & array_obj_ref_1131_word_address_0;
      array_obj_ref_1141_data_0 <= data_out(255 downto 240);
      array_obj_ref_991_data_0 <= data_out(239 downto 224);
      array_obj_ref_1011_data_0 <= data_out(223 downto 208);
      array_obj_ref_1001_data_0 <= data_out(207 downto 192);
      array_obj_ref_1021_data_0 <= data_out(191 downto 176);
      array_obj_ref_1031_data_0 <= data_out(175 downto 160);
      array_obj_ref_1041_data_0 <= data_out(159 downto 144);
      array_obj_ref_1051_data_0 <= data_out(143 downto 128);
      array_obj_ref_1061_data_0 <= data_out(127 downto 112);
      array_obj_ref_1071_data_0 <= data_out(111 downto 96);
      array_obj_ref_1081_data_0 <= data_out(95 downto 80);
      array_obj_ref_1091_data_0 <= data_out(79 downto 64);
      array_obj_ref_1101_data_0 <= data_out(63 downto 48);
      array_obj_ref_1111_data_0 <= data_out(47 downto 32);
      array_obj_ref_1121_data_0 <= data_out(31 downto 16);
      array_obj_ref_1131_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 4,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(3 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 16,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator array_obj_ref_988_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_988_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_load_0:started:   inputs: " & " array_obj_ref_988_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_988_word_address_0));
          --
        end if; 
        if array_obj_ref_988_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_988_load_0:finished:  outputs: " & " array_obj_ref_988_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_988_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1008_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1008_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_load_0:started:   inputs: " & " array_obj_ref_1008_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1008_word_address_0));
          --
        end if; 
        if array_obj_ref_1008_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1008_load_0:finished:  outputs: " & " array_obj_ref_1008_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1008_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_998_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_998_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_load_0:started:   inputs: " & " array_obj_ref_998_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_998_word_address_0));
          --
        end if; 
        if array_obj_ref_998_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_998_load_0:finished:  outputs: " & " array_obj_ref_998_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_998_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1138_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1138_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_load_0:started:   inputs: " & " array_obj_ref_1138_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1138_word_address_0));
          --
        end if; 
        if array_obj_ref_1138_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1138_load_0:finished:  outputs: " & " array_obj_ref_1138_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1138_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1028_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1028_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_load_0:started:   inputs: " & " array_obj_ref_1028_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1028_word_address_0));
          --
        end if; 
        if array_obj_ref_1028_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1028_load_0:finished:  outputs: " & " array_obj_ref_1028_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1028_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1038_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1038_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_load_0:started:   inputs: " & " array_obj_ref_1038_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1038_word_address_0));
          --
        end if; 
        if array_obj_ref_1038_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1038_load_0:finished:  outputs: " & " array_obj_ref_1038_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1038_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1048_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1048_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_load_0:started:   inputs: " & " array_obj_ref_1048_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1048_word_address_0));
          --
        end if; 
        if array_obj_ref_1048_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1048_load_0:finished:  outputs: " & " array_obj_ref_1048_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1048_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1058_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1058_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_load_0:started:   inputs: " & " array_obj_ref_1058_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1058_word_address_0));
          --
        end if; 
        if array_obj_ref_1058_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1058_load_0:finished:  outputs: " & " array_obj_ref_1058_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1058_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1068_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1068_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_load_0:started:   inputs: " & " array_obj_ref_1068_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1068_word_address_0));
          --
        end if; 
        if array_obj_ref_1068_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1068_load_0:finished:  outputs: " & " array_obj_ref_1068_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1068_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1078_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1078_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_load_0:started:   inputs: " & " array_obj_ref_1078_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1078_word_address_0));
          --
        end if; 
        if array_obj_ref_1078_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1078_load_0:finished:  outputs: " & " array_obj_ref_1078_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1078_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1088_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1088_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_load_0:started:   inputs: " & " array_obj_ref_1088_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1088_word_address_0));
          --
        end if; 
        if array_obj_ref_1088_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1088_load_0:finished:  outputs: " & " array_obj_ref_1088_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1088_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1098_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1098_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_load_0:started:   inputs: " & " array_obj_ref_1098_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1098_word_address_0));
          --
        end if; 
        if array_obj_ref_1098_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1098_load_0:finished:  outputs: " & " array_obj_ref_1098_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1098_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1108_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1108_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_load_0:started:   inputs: " & " array_obj_ref_1108_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1108_word_address_0));
          --
        end if; 
        if array_obj_ref_1108_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1108_load_0:finished:  outputs: " & " array_obj_ref_1108_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1108_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1118_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1118_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_load_0:started:   inputs: " & " array_obj_ref_1118_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1118_word_address_0));
          --
        end if; 
        if array_obj_ref_1118_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1118_load_0:finished:  outputs: " & " array_obj_ref_1118_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1118_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1128_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1128_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_load_0:started:   inputs: " & " array_obj_ref_1128_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1128_word_address_0));
          --
        end if; 
        if array_obj_ref_1128_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1128_load_0:finished:  outputs: " & " array_obj_ref_1128_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1128_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (1) : array_obj_ref_988_load_0 array_obj_ref_1008_load_0 array_obj_ref_998_load_0 array_obj_ref_1138_load_0 array_obj_ref_1028_load_0 array_obj_ref_1038_load_0 array_obj_ref_1048_load_0 array_obj_ref_1058_load_0 array_obj_ref_1068_load_0 array_obj_ref_1078_load_0 array_obj_ref_1088_load_0 array_obj_ref_1098_load_0 array_obj_ref_1108_load_0 array_obj_ref_1118_load_0 array_obj_ref_1128_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(59 downto 0);
      signal data_out: std_logic_vector(239 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 14 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 14 downto 0);
      signal guard_vector : std_logic_vector( 14 downto 0);
      constant inBUFs : IntegerArray(14 downto 0) := (14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(14 downto 0) := (14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(14 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false);
      constant guardBuffering: IntegerArray(14 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_988_load_0_req_0,
        array_obj_ref_988_load_0_ack_0,
        array_obj_ref_988_load_0_req_1,
        array_obj_ref_988_load_0_ack_1,
        "array_obj_ref_988_load_0",
        "memory_space_2" ,
        array_obj_ref_988_data_0,
        array_obj_ref_988_word_address_0,
        "array_obj_ref_988_data_0",
        "array_obj_ref_988_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1008_load_0_req_0,
        array_obj_ref_1008_load_0_ack_0,
        array_obj_ref_1008_load_0_req_1,
        array_obj_ref_1008_load_0_ack_1,
        "array_obj_ref_1008_load_0",
        "memory_space_2" ,
        array_obj_ref_1008_data_0,
        array_obj_ref_1008_word_address_0,
        "array_obj_ref_1008_data_0",
        "array_obj_ref_1008_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_998_load_0_req_0,
        array_obj_ref_998_load_0_ack_0,
        array_obj_ref_998_load_0_req_1,
        array_obj_ref_998_load_0_ack_1,
        "array_obj_ref_998_load_0",
        "memory_space_2" ,
        array_obj_ref_998_data_0,
        array_obj_ref_998_word_address_0,
        "array_obj_ref_998_data_0",
        "array_obj_ref_998_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1138_load_0_req_0,
        array_obj_ref_1138_load_0_ack_0,
        array_obj_ref_1138_load_0_req_1,
        array_obj_ref_1138_load_0_ack_1,
        "array_obj_ref_1138_load_0",
        "memory_space_2" ,
        array_obj_ref_1138_data_0,
        array_obj_ref_1138_word_address_0,
        "array_obj_ref_1138_data_0",
        "array_obj_ref_1138_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1028_load_0_req_0,
        array_obj_ref_1028_load_0_ack_0,
        array_obj_ref_1028_load_0_req_1,
        array_obj_ref_1028_load_0_ack_1,
        "array_obj_ref_1028_load_0",
        "memory_space_2" ,
        array_obj_ref_1028_data_0,
        array_obj_ref_1028_word_address_0,
        "array_obj_ref_1028_data_0",
        "array_obj_ref_1028_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1038_load_0_req_0,
        array_obj_ref_1038_load_0_ack_0,
        array_obj_ref_1038_load_0_req_1,
        array_obj_ref_1038_load_0_ack_1,
        "array_obj_ref_1038_load_0",
        "memory_space_2" ,
        array_obj_ref_1038_data_0,
        array_obj_ref_1038_word_address_0,
        "array_obj_ref_1038_data_0",
        "array_obj_ref_1038_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1048_load_0_req_0,
        array_obj_ref_1048_load_0_ack_0,
        array_obj_ref_1048_load_0_req_1,
        array_obj_ref_1048_load_0_ack_1,
        "array_obj_ref_1048_load_0",
        "memory_space_2" ,
        array_obj_ref_1048_data_0,
        array_obj_ref_1048_word_address_0,
        "array_obj_ref_1048_data_0",
        "array_obj_ref_1048_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1058_load_0_req_0,
        array_obj_ref_1058_load_0_ack_0,
        array_obj_ref_1058_load_0_req_1,
        array_obj_ref_1058_load_0_ack_1,
        "array_obj_ref_1058_load_0",
        "memory_space_2" ,
        array_obj_ref_1058_data_0,
        array_obj_ref_1058_word_address_0,
        "array_obj_ref_1058_data_0",
        "array_obj_ref_1058_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1068_load_0_req_0,
        array_obj_ref_1068_load_0_ack_0,
        array_obj_ref_1068_load_0_req_1,
        array_obj_ref_1068_load_0_ack_1,
        "array_obj_ref_1068_load_0",
        "memory_space_2" ,
        array_obj_ref_1068_data_0,
        array_obj_ref_1068_word_address_0,
        "array_obj_ref_1068_data_0",
        "array_obj_ref_1068_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1078_load_0_req_0,
        array_obj_ref_1078_load_0_ack_0,
        array_obj_ref_1078_load_0_req_1,
        array_obj_ref_1078_load_0_ack_1,
        "array_obj_ref_1078_load_0",
        "memory_space_2" ,
        array_obj_ref_1078_data_0,
        array_obj_ref_1078_word_address_0,
        "array_obj_ref_1078_data_0",
        "array_obj_ref_1078_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1088_load_0_req_0,
        array_obj_ref_1088_load_0_ack_0,
        array_obj_ref_1088_load_0_req_1,
        array_obj_ref_1088_load_0_ack_1,
        "array_obj_ref_1088_load_0",
        "memory_space_2" ,
        array_obj_ref_1088_data_0,
        array_obj_ref_1088_word_address_0,
        "array_obj_ref_1088_data_0",
        "array_obj_ref_1088_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1098_load_0_req_0,
        array_obj_ref_1098_load_0_ack_0,
        array_obj_ref_1098_load_0_req_1,
        array_obj_ref_1098_load_0_ack_1,
        "array_obj_ref_1098_load_0",
        "memory_space_2" ,
        array_obj_ref_1098_data_0,
        array_obj_ref_1098_word_address_0,
        "array_obj_ref_1098_data_0",
        "array_obj_ref_1098_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1108_load_0_req_0,
        array_obj_ref_1108_load_0_ack_0,
        array_obj_ref_1108_load_0_req_1,
        array_obj_ref_1108_load_0_ack_1,
        "array_obj_ref_1108_load_0",
        "memory_space_2" ,
        array_obj_ref_1108_data_0,
        array_obj_ref_1108_word_address_0,
        "array_obj_ref_1108_data_0",
        "array_obj_ref_1108_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1118_load_0_req_0,
        array_obj_ref_1118_load_0_ack_0,
        array_obj_ref_1118_load_0_req_1,
        array_obj_ref_1118_load_0_ack_1,
        "array_obj_ref_1118_load_0",
        "memory_space_2" ,
        array_obj_ref_1118_data_0,
        array_obj_ref_1118_word_address_0,
        "array_obj_ref_1118_data_0",
        "array_obj_ref_1118_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1128_load_0_req_0,
        array_obj_ref_1128_load_0_ack_0,
        array_obj_ref_1128_load_0_req_1,
        array_obj_ref_1128_load_0_ack_1,
        "array_obj_ref_1128_load_0",
        "memory_space_2" ,
        array_obj_ref_1128_data_0,
        array_obj_ref_1128_word_address_0,
        "array_obj_ref_1128_data_0",
        "array_obj_ref_1128_word_address_0" -- 
      );
      reqL_unguarded(14) <= array_obj_ref_988_load_0_req_0;
      reqL_unguarded(13) <= array_obj_ref_1008_load_0_req_0;
      reqL_unguarded(12) <= array_obj_ref_998_load_0_req_0;
      reqL_unguarded(11) <= array_obj_ref_1138_load_0_req_0;
      reqL_unguarded(10) <= array_obj_ref_1028_load_0_req_0;
      reqL_unguarded(9) <= array_obj_ref_1038_load_0_req_0;
      reqL_unguarded(8) <= array_obj_ref_1048_load_0_req_0;
      reqL_unguarded(7) <= array_obj_ref_1058_load_0_req_0;
      reqL_unguarded(6) <= array_obj_ref_1068_load_0_req_0;
      reqL_unguarded(5) <= array_obj_ref_1078_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_1088_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1098_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1108_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1118_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1128_load_0_req_0;
      array_obj_ref_988_load_0_ack_0 <= ackL_unguarded(14);
      array_obj_ref_1008_load_0_ack_0 <= ackL_unguarded(13);
      array_obj_ref_998_load_0_ack_0 <= ackL_unguarded(12);
      array_obj_ref_1138_load_0_ack_0 <= ackL_unguarded(11);
      array_obj_ref_1028_load_0_ack_0 <= ackL_unguarded(10);
      array_obj_ref_1038_load_0_ack_0 <= ackL_unguarded(9);
      array_obj_ref_1048_load_0_ack_0 <= ackL_unguarded(8);
      array_obj_ref_1058_load_0_ack_0 <= ackL_unguarded(7);
      array_obj_ref_1068_load_0_ack_0 <= ackL_unguarded(6);
      array_obj_ref_1078_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_1088_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1098_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1108_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1118_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1128_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(14) <= array_obj_ref_988_load_0_req_1;
      reqR_unguarded(13) <= array_obj_ref_1008_load_0_req_1;
      reqR_unguarded(12) <= array_obj_ref_998_load_0_req_1;
      reqR_unguarded(11) <= array_obj_ref_1138_load_0_req_1;
      reqR_unguarded(10) <= array_obj_ref_1028_load_0_req_1;
      reqR_unguarded(9) <= array_obj_ref_1038_load_0_req_1;
      reqR_unguarded(8) <= array_obj_ref_1048_load_0_req_1;
      reqR_unguarded(7) <= array_obj_ref_1058_load_0_req_1;
      reqR_unguarded(6) <= array_obj_ref_1068_load_0_req_1;
      reqR_unguarded(5) <= array_obj_ref_1078_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_1088_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1098_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1108_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1118_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1128_load_0_req_1;
      array_obj_ref_988_load_0_ack_1 <= ackR_unguarded(14);
      array_obj_ref_1008_load_0_ack_1 <= ackR_unguarded(13);
      array_obj_ref_998_load_0_ack_1 <= ackR_unguarded(12);
      array_obj_ref_1138_load_0_ack_1 <= ackR_unguarded(11);
      array_obj_ref_1028_load_0_ack_1 <= ackR_unguarded(10);
      array_obj_ref_1038_load_0_ack_1 <= ackR_unguarded(9);
      array_obj_ref_1048_load_0_ack_1 <= ackR_unguarded(8);
      array_obj_ref_1058_load_0_ack_1 <= ackR_unguarded(7);
      array_obj_ref_1068_load_0_ack_1 <= ackR_unguarded(6);
      array_obj_ref_1078_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_1088_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1098_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1108_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1118_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1128_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_8: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_9: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_10: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_11: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_12: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_13: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_14: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 15, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_988_word_address_0 & array_obj_ref_1008_word_address_0 & array_obj_ref_998_word_address_0 & array_obj_ref_1138_word_address_0 & array_obj_ref_1028_word_address_0 & array_obj_ref_1038_word_address_0 & array_obj_ref_1048_word_address_0 & array_obj_ref_1058_word_address_0 & array_obj_ref_1068_word_address_0 & array_obj_ref_1078_word_address_0 & array_obj_ref_1088_word_address_0 & array_obj_ref_1098_word_address_0 & array_obj_ref_1108_word_address_0 & array_obj_ref_1118_word_address_0 & array_obj_ref_1128_word_address_0;
      array_obj_ref_988_data_0 <= data_out(239 downto 224);
      array_obj_ref_1008_data_0 <= data_out(223 downto 208);
      array_obj_ref_998_data_0 <= data_out(207 downto 192);
      array_obj_ref_1138_data_0 <= data_out(191 downto 176);
      array_obj_ref_1028_data_0 <= data_out(175 downto 160);
      array_obj_ref_1038_data_0 <= data_out(159 downto 144);
      array_obj_ref_1048_data_0 <= data_out(143 downto 128);
      array_obj_ref_1058_data_0 <= data_out(127 downto 112);
      array_obj_ref_1068_data_0 <= data_out(111 downto 96);
      array_obj_ref_1078_data_0 <= data_out(95 downto 80);
      array_obj_ref_1088_data_0 <= data_out(79 downto 64);
      array_obj_ref_1098_data_0 <= data_out(63 downto 48);
      array_obj_ref_1108_data_0 <= data_out(47 downto 32);
      array_obj_ref_1118_data_0 <= data_out(31 downto 16);
      array_obj_ref_1128_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 4,
        num_reqs => 15,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(3 downto 0),
          mtag => memory_space_2_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 15,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logger for split-operator array_obj_ref_1018_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1018_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_load_0:started:   inputs: " & " array_obj_ref_1018_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1018_word_address_0));
          --
        end if; 
        if array_obj_ref_1018_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:mainAcc2:DP:array_obj_ref_1018_load_0:finished:  outputs: " & " array_obj_ref_1018_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1018_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (2) : array_obj_ref_1018_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1018_load_0_req_0,
        array_obj_ref_1018_load_0_ack_0,
        array_obj_ref_1018_load_0_req_1,
        array_obj_ref_1018_load_0_ack_1,
        "array_obj_ref_1018_load_0",
        "memory_space_1" ,
        array_obj_ref_1018_data_0,
        array_obj_ref_1018_word_address_0,
        "array_obj_ref_1018_data_0",
        "array_obj_ref_1018_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_1018_load_0_req_0;
      array_obj_ref_1018_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1018_load_0_req_1;
      array_obj_ref_1018_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1018_word_address_0;
      array_obj_ref_1018_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 4,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(3 downto 0),
          mtag => memory_space_1_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- 
  end Block; -- data_path
  -- 
end mainAcc2_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity memAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    env_mem_request_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    env_mem_request_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    env_mem_request_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    env_mem_response_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    env_mem_response_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    env_mem_response_1_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memAccessDaemon;
architecture memAccessDaemon_arch of memAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal memAccessDaemon_CP_7349_start: Boolean;
  signal memAccessDaemon_CP_7349_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1443_call_req_0 : boolean;
  signal WPIPE_env_mem_response_1_1444_inst_req_0 : boolean;
  signal call_stmt_1443_call_ack_0 : boolean;
  signal do_while_stmt_1417_branch_ack_0 : boolean;
  signal RPIPE_env_mem_request_1_1420_inst_req_1 : boolean;
  signal do_while_stmt_1417_branch_req_0 : boolean;
  signal RPIPE_env_mem_request_1_1420_inst_ack_1 : boolean;
  signal call_stmt_1443_call_req_1 : boolean;
  signal call_stmt_1443_call_ack_1 : boolean;
  signal WPIPE_env_mem_response_1_1444_inst_ack_0 : boolean;
  signal WPIPE_env_mem_response_1_1444_inst_req_1 : boolean;
  signal do_while_stmt_1417_branch_ack_1 : boolean;
  signal WPIPE_env_mem_response_1_1444_inst_ack_1 : boolean;
  signal RPIPE_env_mem_request_1_1420_inst_req_0 : boolean;
  signal RPIPE_env_mem_request_1_1420_inst_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "memAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  memAccessDaemon_CP_7349_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "memAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon_CP_7349_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= memAccessDaemon_CP_7349_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon_CP_7349_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon_CP_7349_start,"memAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon_CP_7349_symbol, "memAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  memAccessDaemon_CP_7349: Block -- control-path 
    signal memAccessDaemon_CP_7349_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    memAccessDaemon_CP_7349_elements(0) <= memAccessDaemon_CP_7349_start;
    memAccessDaemon_CP_7349_symbol <= memAccessDaemon_CP_7349_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1416/do_while_stmt_1417__entry__
      -- CP-element group 0: 	 branch_block_stmt_1416/branch_block_stmt_1416__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1416/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	24 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1416/$exit
      -- CP-element group 1: 	 branch_block_stmt_1416/do_while_stmt_1417__exit__
      -- CP-element group 1: 	 branch_block_stmt_1416/branch_block_stmt_1416__exit__
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(1) <= memAccessDaemon_CP_7349_elements(24);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417__entry__
      -- CP-element group 2: 	 branch_block_stmt_1416/do_while_stmt_1417/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(2) <= memAccessDaemon_CP_7349_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	24 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417__exit__
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_7349_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_back
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_7349_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: 	23 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1416/do_while_stmt_1417/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_exit/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(5) <= memAccessDaemon_CP_7349_elements(21);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	20 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_body_done
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(6) <= memAccessDaemon_CP_7349_elements(20);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(7) <= memAccessDaemon_CP_7349_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(8) <= memAccessDaemon_CP_7349_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon_CP_7349_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Sample/rr
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_env_mem_request_1_1420_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_7382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(10), ack => RPIPE_env_mem_request_1_1420_inst_req_0); -- 
    memAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_7349_elements(9) & memAccessDaemon_CP_7349_elements(13);
      gj_memAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Update/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_env_mem_request_1_1420_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(11), ack => RPIPE_env_mem_request_1_1420_inst_req_1); -- 
    memAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_7349_elements(12) & memAccessDaemon_CP_7349_elements(16);
      gj_memAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Sample/ra
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_env_mem_request_1_1420_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_env_mem_request_1_1420_inst_ack_0, ack => memAccessDaemon_CP_7349_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/RPIPE_env_mem_request_1_1420_update_completed_
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:RPIPE_env_mem_request_1_1420_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_env_mem_request_1_1420_inst_ack_1, ack => memAccessDaemon_CP_7349_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Sample/crr
      -- CP-element group 14: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Sample/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_1443_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(14), ack => call_stmt_1443_call_req_0); -- 
    memAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_7349_elements(13) & memAccessDaemon_CP_7349_elements(16);
      gj_memAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Update/ccr
      -- CP-element group 15: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_update_start_
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_1443_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(15), ack => call_stmt_1443_call_req_1); -- 
    memAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memAccessDaemon_CP_7349_elements(19);
      gj_memAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Sample/cra
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_1443_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1443_call_ack_0, ack => memAccessDaemon_CP_7349_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_Update/cca
      -- CP-element group 17: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/call_stmt_1443_update_completed_
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:call_stmt_1443_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1443_call_ack_1, ack => memAccessDaemon_CP_7349_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Sample/req
      -- CP-element group 18: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_sample_start_
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_env_mem_response_1_1444_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(18), ack => WPIPE_env_mem_response_1_1444_inst_req_0); -- 
    memAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "memAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon_CP_7349_elements(17) & memAccessDaemon_CP_7349_elements(20);
      gj_memAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Update/req
      -- CP-element group 19: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Update/$entry
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_env_mem_response_1_1444_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_env_mem_response_1_1444_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_env_mem_response_1_1444_inst_ack_0, ack => memAccessDaemon_CP_7349_elements(19)); -- 
    req_7415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(19), ack => WPIPE_env_mem_response_1_1444_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (4) 
      -- CP-element group 20: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/$exit
      -- CP-element group 20: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_Update/ack
      -- CP-element group 20: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/WPIPE_env_mem_response_1_1444_update_completed_
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:WPIPE_env_mem_response_1_1444_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_env_mem_response_1_1444_inst_ack_1, ack => memAccessDaemon_CP_7349_elements(20)); -- 
    -- CP-element group 21:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	5 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/loop_body_delay_to_condition_start
      -- CP-element group 21: 	 branch_block_stmt_1416/do_while_stmt_1417/do_while_stmt_1417_loop_body/condition_evaluated
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_1417_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_7373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon_CP_7349_elements(21), ack => do_while_stmt_1417_branch_req_0); -- 
    -- Element group memAccessDaemon_CP_7349_elements(21) is a control-delay.
    cp_element_21_delay: control_delay_element  generic map(name => " 21_delay", delay_value => 1)  port map(req => memAccessDaemon_CP_7349_elements(9), ack => memAccessDaemon_CP_7349_elements(21), clk => clk, reset =>reset);
    -- CP-element group 22:  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_exit/ack
      -- CP-element group 22: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_exit/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_1417_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1417_branch_ack_0, ack => memAccessDaemon_CP_7349_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	5 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_taken/$exit
      -- CP-element group 23: 	 branch_block_stmt_1416/do_while_stmt_1417/loop_taken/ack
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:do_while_stmt_1417_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1417_branch_ack_1, ack => memAccessDaemon_CP_7349_elements(23)); -- 
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	3 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	1 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1416/do_while_stmt_1417/$exit
      -- 
    -- logger for CP element group memAccessDaemon_CP_7349_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon_CP_7349_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon:CP:memAccessDaemon_CP_7349_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon_CP_7349_elements(24) <= memAccessDaemon_CP_7349_elements(3);
    memAccessDaemon_do_while_stmt_1417_terminator_7426: loop_terminator -- 
      generic map (name => " memAccessDaemon_do_while_stmt_1417_terminator_7426", max_iterations_in_flight =>20) 
      port map(loop_body_exit => memAccessDaemon_CP_7349_elements(6),loop_continue => memAccessDaemon_CP_7349_elements(23),loop_terminate => memAccessDaemon_CP_7349_elements(22),loop_back => memAccessDaemon_CP_7349_elements(4),loop_exit => memAccessDaemon_CP_7349_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_7374_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= memAccessDaemon_CP_7349_elements(7);
        preds(1)  <= memAccessDaemon_CP_7349_elements(8);
        entry_tmerge_7374 : transition_merge -- 
          generic map(name => " entry_tmerge_7374")
          port map (preds => preds, symbol_out => memAccessDaemon_CP_7349_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal cmd_1_1421 : std_logic_vector(31 downto 0);
    signal col_index1_1433 : std_logic_vector(4 downto 0);
    signal konst_1448_wire_constant : std_logic_vector(0 downto 0);
    signal rdata1_1443 : std_logic_vector(15 downto 0);
    signal row_index1_1429 : std_logic_vector(5 downto 0);
    signal rwbar1_1437 : std_logic_vector(0 downto 0);
    signal wdata1_1425 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    konst_1448_wire_constant <= "1";
    -- logger for split-operator slice_1424_inst flow-through 
    process(wdata1_1425) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_1424_inst:flowthrough inputs: " & " cmd_1_1421 = "& Convert_SLV_To_Hex_String(cmd_1_1421) & " outputs:" & " wdata1_1425= "  & Convert_SLV_To_Hex_String(wdata1_1425));
      --
    end process; 
    -- flow-through slice operator slice_1424_inst
    wdata1_1425 <= cmd_1_1421(31 downto 16);
    -- logger for split-operator slice_1428_inst flow-through 
    process(row_index1_1429) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_1428_inst:flowthrough inputs: " & " cmd_1_1421 = "& Convert_SLV_To_Hex_String(cmd_1_1421) & " outputs:" & " row_index1_1429= "  & Convert_SLV_To_Hex_String(row_index1_1429));
      --
    end process; 
    -- flow-through slice operator slice_1428_inst
    row_index1_1429 <= cmd_1_1421(15 downto 10);
    -- logger for split-operator slice_1432_inst flow-through 
    process(col_index1_1433) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_1432_inst:flowthrough inputs: " & " cmd_1_1421 = "& Convert_SLV_To_Hex_String(cmd_1_1421) & " outputs:" & " col_index1_1433= "  & Convert_SLV_To_Hex_String(col_index1_1433));
      --
    end process; 
    -- flow-through slice operator slice_1432_inst
    col_index1_1433 <= cmd_1_1421(9 downto 5);
    -- logger for split-operator slice_1436_inst flow-through 
    process(rwbar1_1437) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:slice_1436_inst:flowthrough inputs: " & " cmd_1_1421 = "& Convert_SLV_To_Hex_String(cmd_1_1421) & " outputs:" & " rwbar1_1437= "  & Convert_SLV_To_Hex_String(rwbar1_1437));
      --
    end process; 
    -- flow-through slice operator slice_1436_inst
    rwbar1_1437 <= cmd_1_1421(0 downto 0);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1417_branch_req_0," req0 do_while_stmt_1417_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1417_branch_ack_0," ack0 do_while_stmt_1417_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1417_branch_ack_1," ack1 do_while_stmt_1417_branch");
    do_while_stmt_1417_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1448_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1417_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1417_branch_req_0,
          ack0 => do_while_stmt_1417_branch_ack_0,
          ack1 => do_while_stmt_1417_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_env_mem_request_1_1420_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_env_mem_request_1_1420_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:RPIPE_env_mem_request_1_1420_inst:started:   PipeRead from env_mem_request_1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_env_mem_request_1_1420_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:RPIPE_env_mem_request_1_1420_inst:finished:  outputs: " & " cmd_1_1421= "  & Convert_SLV_To_Hex_String(cmd_1_1421));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_env_mem_request_1_1420_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_env_mem_request_1_1420_inst_req_0;
      RPIPE_env_mem_request_1_1420_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_env_mem_request_1_1420_inst_req_1;
      RPIPE_env_mem_request_1_1420_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_1_1421 <= data_out(31 downto 0);
      env_mem_request_1_read_0_gI: SplitGuardInterface generic map(name => "env_mem_request_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      env_mem_request_1_read_0: InputPortRevised -- 
        generic map ( name => "env_mem_request_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => env_mem_request_1_pipe_read_req(0),
          oack => env_mem_request_1_pipe_read_ack(0),
          odata => env_mem_request_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_env_mem_response_1_1444_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_env_mem_response_1_1444_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:WPIPE_env_mem_response_1_1444_inst:started:   PipeWrite to env_mem_response_1 inputs: " & " rdata1_1443 = "& Convert_SLV_To_Hex_String(rdata1_1443));
          --
        end if; 
        if WPIPE_env_mem_response_1_1444_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:WPIPE_env_mem_response_1_1444_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_env_mem_response_1_1444_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_env_mem_response_1_1444_inst_req_0;
      WPIPE_env_mem_response_1_1444_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_env_mem_response_1_1444_inst_req_1;
      WPIPE_env_mem_response_1_1444_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata1_1443;
      env_mem_response_1_write_0_gI: SplitGuardInterface generic map(name => "env_mem_response_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      env_mem_response_1_write_0: OutputPortRevised -- 
        generic map ( name => "env_mem_response_1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => env_mem_response_1_pipe_write_req(0),
          oack => env_mem_response_1_pipe_write_ack(0),
          odata => env_mem_response_1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_1443_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1443_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:call_stmt_1443_call:started:  Call to module accessMem inputs: " & " rwbar1_1437 = "& Convert_SLV_To_Hex_String(rwbar1_1437) & " row_index1_1429 = "& Convert_SLV_To_Hex_String(row_index1_1429) & " col_index1_1433 = "& Convert_SLV_To_Hex_String(col_index1_1433) & " wdata1_1425 = "& Convert_SLV_To_Hex_String(wdata1_1425));
          --
        end if; 
        if call_stmt_1443_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon:DP:call_stmt_1443_call:finished:  outputs: " & " rdata1_1443= "  & Convert_SLV_To_Hex_String(rdata1_1443));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1443_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1443_call_req_0;
      call_stmt_1443_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1443_call_req_1;
      call_stmt_1443_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar1_1437 & row_index1_1429 & col_index1_1433 & wdata1_1425;
      rdata1_1443 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 28,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 5,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end memAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity memAccessDaemon2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    env_mem_request_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    env_mem_request_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    env_mem_request_2_pipe_read_data : in   std_logic_vector(31 downto 0);
    env_mem_response_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    env_mem_response_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    env_mem_response_2_pipe_write_data : out  std_logic_vector(15 downto 0);
    accessMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessMem_call_acks : in   std_logic_vector(0 downto 0);
    accessMem_call_data : out  std_logic_vector(27 downto 0);
    accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
    accessMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessMem_return_acks : in   std_logic_vector(0 downto 0);
    accessMem_return_data : in   std_logic_vector(15 downto 0);
    accessMem_return_tag :  in   std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memAccessDaemon2;
architecture memAccessDaemon2_arch of memAccessDaemon2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal memAccessDaemon2_CP_7427_start: Boolean;
  signal memAccessDaemon2_CP_7427_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_1453_branch_req_0 : boolean;
  signal call_stmt_1479_call_ack_1 : boolean;
  signal call_stmt_1479_call_req_1 : boolean;
  signal RPIPE_env_mem_request_2_1456_inst_req_0 : boolean;
  signal RPIPE_env_mem_request_2_1456_inst_req_1 : boolean;
  signal RPIPE_env_mem_request_2_1456_inst_ack_1 : boolean;
  signal RPIPE_env_mem_request_2_1456_inst_ack_0 : boolean;
  signal WPIPE_env_mem_response_2_1480_inst_req_0 : boolean;
  signal call_stmt_1479_call_req_0 : boolean;
  signal WPIPE_env_mem_response_2_1480_inst_ack_0 : boolean;
  signal call_stmt_1479_call_ack_0 : boolean;
  signal WPIPE_env_mem_response_2_1480_inst_req_1 : boolean;
  signal WPIPE_env_mem_response_2_1480_inst_ack_1 : boolean;
  signal do_while_stmt_1453_branch_ack_0 : boolean;
  signal do_while_stmt_1453_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "memAccessDaemon2_input_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  memAccessDaemon2_CP_7427_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "memAccessDaemon2_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon2_CP_7427_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= memAccessDaemon2_CP_7427_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memAccessDaemon2_CP_7427_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon2_CP_7427_start,"memAccessDaemon2 cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,memAccessDaemon2_CP_7427_symbol, "memAccessDaemon2 cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  memAccessDaemon2_CP_7427: Block -- control-path 
    signal memAccessDaemon2_CP_7427_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    memAccessDaemon2_CP_7427_elements(0) <= memAccessDaemon2_CP_7427_start;
    memAccessDaemon2_CP_7427_symbol <= memAccessDaemon2_CP_7427_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1452/$entry
      -- CP-element group 0: 	 branch_block_stmt_1452/branch_block_stmt_1452__entry__
      -- CP-element group 0: 	 branch_block_stmt_1452/do_while_stmt_1453__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	24 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1452/$exit
      -- CP-element group 1: 	 branch_block_stmt_1452/branch_block_stmt_1452__exit__
      -- CP-element group 1: 	 branch_block_stmt_1452/do_while_stmt_1453__exit__
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(1) <= memAccessDaemon2_CP_7427_elements(24);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1452/do_while_stmt_1453/$entry
      -- CP-element group 2: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453__entry__
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(2) <= memAccessDaemon2_CP_7427_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	24 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453__exit__
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon2_CP_7427_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_back
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon2_CP_7427_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	21 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: 	23 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1452/do_while_stmt_1453/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_taken/$entry
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(5) <= memAccessDaemon2_CP_7427_elements(21);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	20 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_body_done
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(6) <= memAccessDaemon2_CP_7427_elements(20);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(7) <= memAccessDaemon2_CP_7427_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(8) <= memAccessDaemon2_CP_7427_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/$entry
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memAccessDaemon2_CP_7427_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_sample_start_
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:RPIPE_env_mem_request_2_1456_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_7460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(10), ack => RPIPE_env_mem_request_2_1456_inst_req_0); -- 
    memAccessDaemon2_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 20,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "memAccessDaemon2_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon2_CP_7427_elements(9) & memAccessDaemon2_CP_7427_elements(13);
      gj_memAccessDaemon2_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Update/cr
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:RPIPE_env_mem_request_2_1456_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_7465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(11), ack => RPIPE_env_mem_request_2_1456_inst_req_1); -- 
    memAccessDaemon2_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "memAccessDaemon2_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon2_CP_7427_elements(12) & memAccessDaemon2_CP_7427_elements(16);
      gj_memAccessDaemon2_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Sample/ra
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:RPIPE_env_mem_request_2_1456_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_7461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_env_mem_request_2_1456_inst_ack_0, ack => memAccessDaemon2_CP_7427_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/RPIPE_env_mem_request_2_1456_Update/ca
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:RPIPE_env_mem_request_2_1456_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_7466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_env_mem_request_2_1456_inst_ack_1, ack => memAccessDaemon2_CP_7427_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Sample/crr
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:call_stmt_1479_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_7474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_7474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(14), ack => call_stmt_1479_call_req_0); -- 
    memAccessDaemon2_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "memAccessDaemon2_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon2_CP_7427_elements(13) & memAccessDaemon2_CP_7427_elements(16);
      gj_memAccessDaemon2_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Update/ccr
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:call_stmt_1479_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_7479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_7479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(15), ack => call_stmt_1479_call_req_1); -- 
    memAccessDaemon2_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "memAccessDaemon2_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memAccessDaemon2_CP_7427_elements(19);
      gj_memAccessDaemon2_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Sample/cra
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:call_stmt_1479_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_7475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1479_call_ack_0, ack => memAccessDaemon2_CP_7427_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Update/cca
      -- CP-element group 17: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/call_stmt_1479_update_completed_
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:call_stmt_1479_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_7480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1479_call_ack_1, ack => memAccessDaemon2_CP_7427_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Sample/req
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:WPIPE_env_mem_response_2_1480_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_7488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(18), ack => WPIPE_env_mem_response_2_1480_inst_req_0); -- 
    memAccessDaemon2_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "memAccessDaemon2_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memAccessDaemon2_CP_7427_elements(17) & memAccessDaemon2_CP_7427_elements(20);
      gj_memAccessDaemon2_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Sample/ack
      -- CP-element group 19: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Update/req
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:WPIPE_env_mem_response_2_1480_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:WPIPE_env_mem_response_2_1480_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_env_mem_response_2_1480_inst_ack_0, ack => memAccessDaemon2_CP_7427_elements(19)); -- 
    req_7493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(19), ack => WPIPE_env_mem_response_2_1480_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (4) 
      -- CP-element group 20: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/$exit
      -- CP-element group 20: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/WPIPE_env_mem_response_2_1480_Update/ack
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:WPIPE_env_mem_response_2_1480_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_env_mem_response_2_1480_inst_ack_1, ack => memAccessDaemon2_CP_7427_elements(20)); -- 
    -- CP-element group 21:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	5 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/condition_evaluated
      -- CP-element group 21: 	 branch_block_stmt_1452/do_while_stmt_1453/do_while_stmt_1453_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:do_while_stmt_1453_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_7451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_7451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memAccessDaemon2_CP_7427_elements(21), ack => do_while_stmt_1453_branch_req_0); -- 
    -- Element group memAccessDaemon2_CP_7427_elements(21) is a control-delay.
    cp_element_21_delay: control_delay_element  generic map(name => " 21_delay", delay_value => 1)  port map(req => memAccessDaemon2_CP_7427_elements(9), ack => memAccessDaemon2_CP_7427_elements(21), clk => clk, reset =>reset);
    -- CP-element group 22:  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	5 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_exit/$exit
      -- CP-element group 22: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_exit/ack
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:do_while_stmt_1453_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_7499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1453_branch_ack_0, ack => memAccessDaemon2_CP_7427_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	5 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_taken/$exit
      -- CP-element group 23: 	 branch_block_stmt_1452/do_while_stmt_1453/loop_taken/ack
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:do_while_stmt_1453_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_7503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1453_branch_ack_1, ack => memAccessDaemon2_CP_7427_elements(23)); -- 
    -- CP-element group 24:  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	3 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	1 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1452/do_while_stmt_1453/$exit
      -- 
    -- logger for CP element group memAccessDaemon2_CP_7427_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memAccessDaemon2_CP_7427_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memAccessDaemon2:CP:memAccessDaemon2_CP_7427_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    memAccessDaemon2_CP_7427_elements(24) <= memAccessDaemon2_CP_7427_elements(3);
    memAccessDaemon2_do_while_stmt_1453_terminator_7504: loop_terminator -- 
      generic map (name => " memAccessDaemon2_do_while_stmt_1453_terminator_7504", max_iterations_in_flight =>20) 
      port map(loop_body_exit => memAccessDaemon2_CP_7427_elements(6),loop_continue => memAccessDaemon2_CP_7427_elements(23),loop_terminate => memAccessDaemon2_CP_7427_elements(22),loop_back => memAccessDaemon2_CP_7427_elements(4),loop_exit => memAccessDaemon2_CP_7427_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_7452_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= memAccessDaemon2_CP_7427_elements(7);
        preds(1)  <= memAccessDaemon2_CP_7427_elements(8);
        entry_tmerge_7452 : transition_merge -- 
          generic map(name => " entry_tmerge_7452")
          port map (preds => preds, symbol_out => memAccessDaemon2_CP_7427_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal cmd_2_1457 : std_logic_vector(31 downto 0);
    signal col_index2_1469 : std_logic_vector(4 downto 0);
    signal konst_1484_wire_constant : std_logic_vector(0 downto 0);
    signal rdata2_1479 : std_logic_vector(15 downto 0);
    signal row_index2_1465 : std_logic_vector(5 downto 0);
    signal rwbar2_1473 : std_logic_vector(0 downto 0);
    signal wdata2_1461 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    konst_1484_wire_constant <= "1";
    -- logger for split-operator slice_1460_inst flow-through 
    process(wdata2_1461) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:slice_1460_inst:flowthrough inputs: " & " cmd_2_1457 = "& Convert_SLV_To_Hex_String(cmd_2_1457) & " outputs:" & " wdata2_1461= "  & Convert_SLV_To_Hex_String(wdata2_1461));
      --
    end process; 
    -- flow-through slice operator slice_1460_inst
    wdata2_1461 <= cmd_2_1457(31 downto 16);
    -- logger for split-operator slice_1464_inst flow-through 
    process(row_index2_1465) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:slice_1464_inst:flowthrough inputs: " & " cmd_2_1457 = "& Convert_SLV_To_Hex_String(cmd_2_1457) & " outputs:" & " row_index2_1465= "  & Convert_SLV_To_Hex_String(row_index2_1465));
      --
    end process; 
    -- flow-through slice operator slice_1464_inst
    row_index2_1465 <= cmd_2_1457(15 downto 10);
    -- logger for split-operator slice_1468_inst flow-through 
    process(col_index2_1469) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:slice_1468_inst:flowthrough inputs: " & " cmd_2_1457 = "& Convert_SLV_To_Hex_String(cmd_2_1457) & " outputs:" & " col_index2_1469= "  & Convert_SLV_To_Hex_String(col_index2_1469));
      --
    end process; 
    -- flow-through slice operator slice_1468_inst
    col_index2_1469 <= cmd_2_1457(9 downto 5);
    -- logger for split-operator slice_1472_inst flow-through 
    process(rwbar2_1473) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:slice_1472_inst:flowthrough inputs: " & " cmd_2_1457 = "& Convert_SLV_To_Hex_String(cmd_2_1457) & " outputs:" & " rwbar2_1473= "  & Convert_SLV_To_Hex_String(rwbar2_1473));
      --
    end process; 
    -- flow-through slice operator slice_1472_inst
    rwbar2_1473 <= cmd_2_1457(0 downto 0);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1453_branch_req_0," req0 do_while_stmt_1453_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1453_branch_ack_0," ack0 do_while_stmt_1453_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1453_branch_ack_1," ack1 do_while_stmt_1453_branch");
    do_while_stmt_1453_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1484_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1453_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1453_branch_req_0,
          ack0 => do_while_stmt_1453_branch_ack_0,
          ack1 => do_while_stmt_1453_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_env_mem_request_2_1456_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_env_mem_request_2_1456_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:RPIPE_env_mem_request_2_1456_inst:started:   PipeRead from env_mem_request_2 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_env_mem_request_2_1456_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:RPIPE_env_mem_request_2_1456_inst:finished:  outputs: " & " cmd_2_1457= "  & Convert_SLV_To_Hex_String(cmd_2_1457));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_env_mem_request_2_1456_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_env_mem_request_2_1456_inst_req_0;
      RPIPE_env_mem_request_2_1456_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_env_mem_request_2_1456_inst_req_1;
      RPIPE_env_mem_request_2_1456_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      cmd_2_1457 <= data_out(31 downto 0);
      env_mem_request_2_read_0_gI: SplitGuardInterface generic map(name => "env_mem_request_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      env_mem_request_2_read_0: InputPortRevised -- 
        generic map ( name => "env_mem_request_2_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => env_mem_request_2_pipe_read_req(0),
          oack => env_mem_request_2_pipe_read_ack(0),
          odata => env_mem_request_2_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_env_mem_response_2_1480_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_env_mem_response_2_1480_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:WPIPE_env_mem_response_2_1480_inst:started:   PipeWrite to env_mem_response_2 inputs: " & " rdata2_1479 = "& Convert_SLV_To_Hex_String(rdata2_1479));
          --
        end if; 
        if WPIPE_env_mem_response_2_1480_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:WPIPE_env_mem_response_2_1480_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_env_mem_response_2_1480_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_env_mem_response_2_1480_inst_req_0;
      WPIPE_env_mem_response_2_1480_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_env_mem_response_2_1480_inst_req_1;
      WPIPE_env_mem_response_2_1480_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= rdata2_1479;
      env_mem_response_2_write_0_gI: SplitGuardInterface generic map(name => "env_mem_response_2_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      env_mem_response_2_write_0: OutputPortRevised -- 
        generic map ( name => "env_mem_response_2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => env_mem_response_2_pipe_write_req(0),
          oack => env_mem_response_2_pipe_write_ack(0),
          odata => env_mem_response_2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_1479_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1479_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:call_stmt_1479_call:started:  Call to module accessMem inputs: " & " rwbar2_1473 = "& Convert_SLV_To_Hex_String(rwbar2_1473) & " row_index2_1465 = "& Convert_SLV_To_Hex_String(row_index2_1465) & " col_index2_1469 = "& Convert_SLV_To_Hex_String(col_index2_1469) & " wdata2_1461 = "& Convert_SLV_To_Hex_String(wdata2_1461));
          --
        end if; 
        if call_stmt_1479_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memAccessDaemon2:DP:call_stmt_1479_call:finished:  outputs: " & " rdata2_1479= "  & Convert_SLV_To_Hex_String(rdata2_1479));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1479_call 
    accessMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 7);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1479_call_req_0;
      call_stmt_1479_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1479_call_req_1;
      call_stmt_1479_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rwbar2_1473 & row_index2_1465 & col_index2_1469 & wdata2_1461;
      rdata2_1479 <= data_out(15 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 28,
        owidth => 28,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 5,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMem_call_reqs(0),
          ackR => accessMem_call_acks(0),
          dataR => accessMem_call_data(27 downto 0),
          tagR => accessMem_call_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 5,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMem_return_acks(0), -- cross-over
          ackL => accessMem_return_reqs(0), -- cross-over
          dataL => accessMem_return_data(15 downto 0),
          tagL => accessMem_return_tag(4 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end memAccessDaemon2_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    acc_mem_request_1_pipe_write_data: in std_logic_vector(31 downto 0);
    acc_mem_request_1_pipe_write_req : in std_logic_vector(0 downto 0);
    acc_mem_request_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    acc_mem_response_1_pipe_read_data: out std_logic_vector(15 downto 0);
    acc_mem_response_1_pipe_read_req : in std_logic_vector(0 downto 0);
    acc_mem_response_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    accelerator_done_pipe_read_data: out std_logic_vector(15 downto 0);
    accelerator_done_pipe_read_req : in std_logic_vector(0 downto 0);
    accelerator_done_pipe_read_ack : out std_logic_vector(0 downto 0);
    env_mem_request_1_pipe_write_data: in std_logic_vector(31 downto 0);
    env_mem_request_1_pipe_write_req : in std_logic_vector(0 downto 0);
    env_mem_request_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    env_mem_request_2_pipe_write_data: in std_logic_vector(31 downto 0);
    env_mem_request_2_pipe_write_req : in std_logic_vector(0 downto 0);
    env_mem_request_2_pipe_write_ack : out std_logic_vector(0 downto 0);
    env_mem_response_1_pipe_read_data: out std_logic_vector(15 downto 0);
    env_mem_response_1_pipe_read_req : in std_logic_vector(0 downto 0);
    env_mem_response_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    env_mem_response_2_pipe_read_data: out std_logic_vector(15 downto 0);
    env_mem_response_2_pipe_read_req : in std_logic_vector(0 downto 0);
    env_mem_response_2_pipe_read_ack : out std_logic_vector(0 downto 0);
    read_sums_pipe_read_data: out std_logic_vector(15 downto 0);
    read_sums_pipe_read_req : in std_logic_vector(0 downto 0);
    read_sums_pipe_read_ack : out std_logic_vector(0 downto 0);
    start_accelerator_pipe_write_data: in std_logic_vector(15 downto 0);
    start_accelerator_pipe_write_req : in std_logic_vector(0 downto 0);
    start_accelerator_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(7 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(7 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(43 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(15 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module accMemAccessDaemon
  component accMemAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      acc_mem_request_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      acc_mem_request_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      acc_mem_request_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      acc_mem_response_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      acc_mem_response_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      acc_mem_response_1_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accMemAccessDaemon
  signal accMemAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accMemAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal accMemAccessDaemon_start_req : std_logic;
  signal accMemAccessDaemon_start_ack : std_logic;
  signal accMemAccessDaemon_fin_req   : std_logic;
  signal accMemAccessDaemon_fin_ack : std_logic;
  -- declarations related to module accelerator
  component accelerator is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_accelerator_pipe_read_req : out  std_logic_vector(0 downto 0);
      start_accelerator_pipe_read_ack : in   std_logic_vector(0 downto 0);
      start_accelerator_pipe_read_data : in   std_logic_vector(15 downto 0);
      accelerator_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      accelerator_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      accelerator_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      read_sums_pipe_write_req : out  std_logic_vector(0 downto 0);
      read_sums_pipe_write_ack : in   std_logic_vector(0 downto 0);
      read_sums_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      initIfMaps_call_reqs : out  std_logic_vector(0 downto 0);
      initIfMaps_call_acks : in   std_logic_vector(0 downto 0);
      initIfMaps_call_data : out  std_logic_vector(13 downto 0);
      initIfMaps_call_tag  :  out  std_logic_vector(0 downto 0);
      initIfMaps_return_reqs : out  std_logic_vector(0 downto 0);
      initIfMaps_return_acks : in   std_logic_vector(0 downto 0);
      initIfMaps_return_data : in   std_logic_vector(1 downto 0);
      initIfMaps_return_tag :  in   std_logic_vector(0 downto 0);
      initFilter_call_reqs : out  std_logic_vector(0 downto 0);
      initFilter_call_acks : in   std_logic_vector(0 downto 0);
      initFilter_call_data : out  std_logic_vector(5 downto 0);
      initFilter_call_tag  :  out  std_logic_vector(0 downto 0);
      initFilter_return_reqs : out  std_logic_vector(0 downto 0);
      initFilter_return_acks : in   std_logic_vector(0 downto 0);
      initFilter_return_data : in   std_logic_vector(1 downto 0);
      initFilter_return_tag :  in   std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_call_reqs : out  std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_call_acks : in   std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_call_data : out  std_logic_vector(6 downto 0);
      cal_col_to_be_replaced_call_tag  :  out  std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_return_reqs : out  std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_return_acks : in   std_logic_vector(0 downto 0);
      cal_col_to_be_replaced_return_data : in   std_logic_vector(1 downto 0);
      cal_col_to_be_replaced_return_tag :  in   std_logic_vector(0 downto 0);
      mainAcc_call_reqs : out  std_logic_vector(0 downto 0);
      mainAcc_call_acks : in   std_logic_vector(0 downto 0);
      mainAcc_call_data : out  std_logic_vector(12 downto 0);
      mainAcc_call_tag  :  out  std_logic_vector(0 downto 0);
      mainAcc_return_reqs : out  std_logic_vector(0 downto 0);
      mainAcc_return_acks : in   std_logic_vector(0 downto 0);
      mainAcc_return_data : in   std_logic_vector(15 downto 0);
      mainAcc_return_tag :  in   std_logic_vector(0 downto 0);
      mainAcc2_call_reqs : out  std_logic_vector(0 downto 0);
      mainAcc2_call_acks : in   std_logic_vector(0 downto 0);
      mainAcc2_call_data : out  std_logic_vector(12 downto 0);
      mainAcc2_call_tag  :  out  std_logic_vector(0 downto 0);
      mainAcc2_return_reqs : out  std_logic_vector(0 downto 0);
      mainAcc2_return_acks : in   std_logic_vector(0 downto 0);
      mainAcc2_return_data : in   std_logic_vector(15 downto 0);
      mainAcc2_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accelerator
  signal accelerator_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accelerator_tag_out   : std_logic_vector(1 downto 0);
  signal accelerator_start_req : std_logic;
  signal accelerator_start_ack : std_logic;
  signal accelerator_fin_req   : std_logic;
  signal accelerator_fin_ack : std_logic;
  -- declarations related to module accessMem
  component accessMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      read_write_bar_1 : in  std_logic_vector(0 downto 0);
      row_index : in  std_logic_vector(5 downto 0);
      col_index : in  std_logic_vector(4 downto 0);
      write_data_1 : in  std_logic_vector(15 downto 0);
      read_data_1 : out  std_logic_vector(15 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMem
  signal accessMem_read_write_bar_1 :  std_logic_vector(0 downto 0);
  signal accessMem_row_index :  std_logic_vector(5 downto 0);
  signal accessMem_col_index :  std_logic_vector(4 downto 0);
  signal accessMem_write_data_1 :  std_logic_vector(15 downto 0);
  signal accessMem_read_data_1 :  std_logic_vector(15 downto 0);
  signal accessMem_in_args    : std_logic_vector(27 downto 0);
  signal accessMem_out_args   : std_logic_vector(15 downto 0);
  signal accessMem_tag_in    : std_logic_vector(7 downto 0) := (others => '0');
  signal accessMem_tag_out   : std_logic_vector(7 downto 0);
  signal accessMem_start_req : std_logic;
  signal accessMem_start_ack : std_logic;
  signal accessMem_fin_req   : std_logic;
  signal accessMem_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMem
  signal accessMem_call_reqs: std_logic_vector(5 downto 0);
  signal accessMem_call_acks: std_logic_vector(5 downto 0);
  signal accessMem_return_reqs: std_logic_vector(5 downto 0);
  signal accessMem_return_acks: std_logic_vector(5 downto 0);
  signal accessMem_call_data: std_logic_vector(167 downto 0);
  signal accessMem_call_tag: std_logic_vector(29 downto 0);
  signal accessMem_return_data: std_logic_vector(95 downto 0);
  signal accessMem_return_tag: std_logic_vector(29 downto 0);
  -- declarations related to module cal_col_to_be_replaced
  component cal_col_to_be_replaced is -- 
    generic (tag_length : integer); 
    port ( -- 
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      new_col_to_be_replaced : out  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module cal_col_to_be_replaced
  signal cal_col_to_be_replaced_J :  std_logic_vector(4 downto 0);
  signal cal_col_to_be_replaced_col_to_be_replaced :  std_logic_vector(1 downto 0);
  signal cal_col_to_be_replaced_new_col_to_be_replaced :  std_logic_vector(1 downto 0);
  signal cal_col_to_be_replaced_in_args    : std_logic_vector(6 downto 0);
  signal cal_col_to_be_replaced_out_args   : std_logic_vector(1 downto 0);
  signal cal_col_to_be_replaced_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal cal_col_to_be_replaced_tag_out   : std_logic_vector(1 downto 0);
  signal cal_col_to_be_replaced_start_req : std_logic;
  signal cal_col_to_be_replaced_start_ack : std_logic;
  signal cal_col_to_be_replaced_fin_req   : std_logic;
  signal cal_col_to_be_replaced_fin_ack : std_logic;
  -- caller side aggregated signals for module cal_col_to_be_replaced
  signal cal_col_to_be_replaced_call_reqs: std_logic_vector(0 downto 0);
  signal cal_col_to_be_replaced_call_acks: std_logic_vector(0 downto 0);
  signal cal_col_to_be_replaced_return_reqs: std_logic_vector(0 downto 0);
  signal cal_col_to_be_replaced_return_acks: std_logic_vector(0 downto 0);
  signal cal_col_to_be_replaced_call_data: std_logic_vector(6 downto 0);
  signal cal_col_to_be_replaced_call_tag: std_logic_vector(0 downto 0);
  signal cal_col_to_be_replaced_return_data: std_logic_vector(1 downto 0);
  signal cal_col_to_be_replaced_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module initFilter
  component initFilter is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_row_filter : in  std_logic_vector(5 downto 0);
      filter_initialized : out  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initFilter
  signal initFilter_start_row_filter :  std_logic_vector(5 downto 0);
  signal initFilter_filter_initialized :  std_logic_vector(1 downto 0);
  signal initFilter_in_args    : std_logic_vector(5 downto 0);
  signal initFilter_out_args   : std_logic_vector(1 downto 0);
  signal initFilter_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initFilter_tag_out   : std_logic_vector(1 downto 0);
  signal initFilter_start_req : std_logic;
  signal initFilter_start_ack : std_logic;
  signal initFilter_fin_req   : std_logic;
  signal initFilter_fin_ack : std_logic;
  -- caller side aggregated signals for module initFilter
  signal initFilter_call_reqs: std_logic_vector(0 downto 0);
  signal initFilter_call_acks: std_logic_vector(0 downto 0);
  signal initFilter_return_reqs: std_logic_vector(0 downto 0);
  signal initFilter_return_acks: std_logic_vector(0 downto 0);
  signal initFilter_call_data: std_logic_vector(5 downto 0);
  signal initFilter_call_tag: std_logic_vector(0 downto 0);
  signal initFilter_return_data: std_logic_vector(1 downto 0);
  signal initFilter_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module initIfMaps
  component initIfMaps is -- 
    generic (tag_length : integer); 
    port ( -- 
      start : in  std_logic_vector(0 downto 0);
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      finished : out  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module initIfMaps
  signal initIfMaps_start :  std_logic_vector(0 downto 0);
  signal initIfMaps_I :  std_logic_vector(5 downto 0);
  signal initIfMaps_J :  std_logic_vector(4 downto 0);
  signal initIfMaps_col_to_be_replaced :  std_logic_vector(1 downto 0);
  signal initIfMaps_finished :  std_logic_vector(1 downto 0);
  signal initIfMaps_in_args    : std_logic_vector(13 downto 0);
  signal initIfMaps_out_args   : std_logic_vector(1 downto 0);
  signal initIfMaps_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal initIfMaps_tag_out   : std_logic_vector(1 downto 0);
  signal initIfMaps_start_req : std_logic;
  signal initIfMaps_start_ack : std_logic;
  signal initIfMaps_fin_req   : std_logic;
  signal initIfMaps_fin_ack : std_logic;
  -- caller side aggregated signals for module initIfMaps
  signal initIfMaps_call_reqs: std_logic_vector(0 downto 0);
  signal initIfMaps_call_acks: std_logic_vector(0 downto 0);
  signal initIfMaps_return_reqs: std_logic_vector(0 downto 0);
  signal initIfMaps_return_acks: std_logic_vector(0 downto 0);
  signal initIfMaps_call_data: std_logic_vector(13 downto 0);
  signal initIfMaps_call_tag: std_logic_vector(0 downto 0);
  signal initIfMaps_return_data: std_logic_vector(1 downto 0);
  signal initIfMaps_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module mainAcc
  component mainAcc is -- 
    generic (tag_length : integer); 
    port ( -- 
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      ofmap_pixel : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module mainAcc
  signal mainAcc_I :  std_logic_vector(5 downto 0);
  signal mainAcc_J :  std_logic_vector(4 downto 0);
  signal mainAcc_col_to_be_replaced :  std_logic_vector(1 downto 0);
  signal mainAcc_ofmap_pixel :  std_logic_vector(15 downto 0);
  signal mainAcc_in_args    : std_logic_vector(12 downto 0);
  signal mainAcc_out_args   : std_logic_vector(15 downto 0);
  signal mainAcc_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal mainAcc_tag_out   : std_logic_vector(1 downto 0);
  signal mainAcc_start_req : std_logic;
  signal mainAcc_start_ack : std_logic;
  signal mainAcc_fin_req   : std_logic;
  signal mainAcc_fin_ack : std_logic;
  -- caller side aggregated signals for module mainAcc
  signal mainAcc_call_reqs: std_logic_vector(0 downto 0);
  signal mainAcc_call_acks: std_logic_vector(0 downto 0);
  signal mainAcc_return_reqs: std_logic_vector(0 downto 0);
  signal mainAcc_return_acks: std_logic_vector(0 downto 0);
  signal mainAcc_call_data: std_logic_vector(12 downto 0);
  signal mainAcc_call_tag: std_logic_vector(0 downto 0);
  signal mainAcc_return_data: std_logic_vector(15 downto 0);
  signal mainAcc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module mainAcc2
  component mainAcc2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      I : in  std_logic_vector(5 downto 0);
      J : in  std_logic_vector(4 downto 0);
      col_to_be_replaced : in  std_logic_vector(1 downto 0);
      ofmap_pixel : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(3 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module mainAcc2
  signal mainAcc2_I :  std_logic_vector(5 downto 0);
  signal mainAcc2_J :  std_logic_vector(4 downto 0);
  signal mainAcc2_col_to_be_replaced :  std_logic_vector(1 downto 0);
  signal mainAcc2_ofmap_pixel :  std_logic_vector(15 downto 0);
  signal mainAcc2_in_args    : std_logic_vector(12 downto 0);
  signal mainAcc2_out_args   : std_logic_vector(15 downto 0);
  signal mainAcc2_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal mainAcc2_tag_out   : std_logic_vector(1 downto 0);
  signal mainAcc2_start_req : std_logic;
  signal mainAcc2_start_ack : std_logic;
  signal mainAcc2_fin_req   : std_logic;
  signal mainAcc2_fin_ack : std_logic;
  -- caller side aggregated signals for module mainAcc2
  signal mainAcc2_call_reqs: std_logic_vector(0 downto 0);
  signal mainAcc2_call_acks: std_logic_vector(0 downto 0);
  signal mainAcc2_return_reqs: std_logic_vector(0 downto 0);
  signal mainAcc2_return_acks: std_logic_vector(0 downto 0);
  signal mainAcc2_call_data: std_logic_vector(12 downto 0);
  signal mainAcc2_call_tag: std_logic_vector(0 downto 0);
  signal mainAcc2_return_data: std_logic_vector(15 downto 0);
  signal mainAcc2_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module memAccessDaemon
  component memAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      env_mem_request_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      env_mem_request_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      env_mem_request_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      env_mem_response_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      env_mem_response_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      env_mem_response_1_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module memAccessDaemon
  signal memAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal memAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal memAccessDaemon_start_req : std_logic;
  signal memAccessDaemon_start_ack : std_logic;
  signal memAccessDaemon_fin_req   : std_logic;
  signal memAccessDaemon_fin_ack : std_logic;
  -- declarations related to module memAccessDaemon2
  component memAccessDaemon2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      env_mem_request_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      env_mem_request_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      env_mem_request_2_pipe_read_data : in   std_logic_vector(31 downto 0);
      env_mem_response_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      env_mem_response_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      env_mem_response_2_pipe_write_data : out  std_logic_vector(15 downto 0);
      accessMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessMem_call_acks : in   std_logic_vector(0 downto 0);
      accessMem_call_data : out  std_logic_vector(27 downto 0);
      accessMem_call_tag  :  out  std_logic_vector(4 downto 0);
      accessMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessMem_return_acks : in   std_logic_vector(0 downto 0);
      accessMem_return_data : in   std_logic_vector(15 downto 0);
      accessMem_return_tag :  in   std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module memAccessDaemon2
  signal memAccessDaemon2_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal memAccessDaemon2_tag_out   : std_logic_vector(1 downto 0);
  signal memAccessDaemon2_start_req : std_logic;
  signal memAccessDaemon2_start_ack : std_logic;
  signal memAccessDaemon2_fin_req   : std_logic;
  signal memAccessDaemon2_fin_ack : std_logic;
  -- aggregate signals for read from pipe acc_mem_request_1
  signal acc_mem_request_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal acc_mem_request_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal acc_mem_request_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe acc_mem_response_1
  signal acc_mem_response_1_pipe_write_data: std_logic_vector(15 downto 0);
  signal acc_mem_response_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal acc_mem_response_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe accelerator_done
  signal accelerator_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal accelerator_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal accelerator_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe env_mem_request_1
  signal env_mem_request_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal env_mem_request_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal env_mem_request_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe env_mem_request_2
  signal env_mem_request_2_pipe_read_data: std_logic_vector(31 downto 0);
  signal env_mem_request_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal env_mem_request_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe env_mem_response_1
  signal env_mem_response_1_pipe_write_data: std_logic_vector(15 downto 0);
  signal env_mem_response_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal env_mem_response_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe env_mem_response_2
  signal env_mem_response_2_pipe_write_data: std_logic_vector(15 downto 0);
  signal env_mem_response_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal env_mem_response_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe read_sums
  signal read_sums_pipe_write_data: std_logic_vector(15 downto 0);
  signal read_sums_pipe_write_req: std_logic_vector(0 downto 0);
  signal read_sums_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe start_accelerator
  signal start_accelerator_pipe_read_data: std_logic_vector(15 downto 0);
  signal start_accelerator_pipe_read_req: std_logic_vector(0 downto 0);
  signal start_accelerator_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module accMemAccessDaemon
  accMemAccessDaemon_instance:accMemAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => accMemAccessDaemon_start_req,
      start_ack => accMemAccessDaemon_start_ack,
      fin_req => accMemAccessDaemon_fin_req,
      fin_ack => accMemAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      acc_mem_request_1_pipe_read_req => acc_mem_request_1_pipe_read_req(0 downto 0),
      acc_mem_request_1_pipe_read_ack => acc_mem_request_1_pipe_read_ack(0 downto 0),
      acc_mem_request_1_pipe_read_data => acc_mem_request_1_pipe_read_data(31 downto 0),
      acc_mem_response_1_pipe_write_req => acc_mem_response_1_pipe_write_req(0 downto 0),
      acc_mem_response_1_pipe_write_ack => acc_mem_response_1_pipe_write_ack(0 downto 0),
      acc_mem_response_1_pipe_write_data => acc_mem_response_1_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(5 downto 5),
      accessMem_call_acks => accessMem_call_acks(5 downto 5),
      accessMem_call_data => accessMem_call_data(167 downto 140),
      accessMem_call_tag => accessMem_call_tag(29 downto 25),
      accessMem_return_reqs => accessMem_return_reqs(5 downto 5),
      accessMem_return_acks => accessMem_return_acks(5 downto 5),
      accessMem_return_data => accessMem_return_data(95 downto 80),
      accessMem_return_tag => accessMem_return_tag(29 downto 25),
      tag_in => accMemAccessDaemon_tag_in,
      tag_out => accMemAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  accMemAccessDaemon_tag_in <= (others => '0');
  accMemAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => accMemAccessDaemon_start_req, start_ack => accMemAccessDaemon_start_ack,  fin_req => accMemAccessDaemon_fin_req,  fin_ack => accMemAccessDaemon_fin_ack);
  -- module accelerator
  accelerator_instance:accelerator-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => accelerator_start_req,
      start_ack => accelerator_start_ack,
      fin_req => accelerator_fin_req,
      fin_ack => accelerator_fin_ack,
      clk => clk,
      reset => reset,
      start_accelerator_pipe_read_req => start_accelerator_pipe_read_req(0 downto 0),
      start_accelerator_pipe_read_ack => start_accelerator_pipe_read_ack(0 downto 0),
      start_accelerator_pipe_read_data => start_accelerator_pipe_read_data(15 downto 0),
      accelerator_done_pipe_write_req => accelerator_done_pipe_write_req(0 downto 0),
      accelerator_done_pipe_write_ack => accelerator_done_pipe_write_ack(0 downto 0),
      accelerator_done_pipe_write_data => accelerator_done_pipe_write_data(15 downto 0),
      read_sums_pipe_write_req => read_sums_pipe_write_req(0 downto 0),
      read_sums_pipe_write_ack => read_sums_pipe_write_ack(0 downto 0),
      read_sums_pipe_write_data => read_sums_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(0 downto 0),
      accessMem_call_acks => accessMem_call_acks(0 downto 0),
      accessMem_call_data => accessMem_call_data(27 downto 0),
      accessMem_call_tag => accessMem_call_tag(4 downto 0),
      accessMem_return_reqs => accessMem_return_reqs(0 downto 0),
      accessMem_return_acks => accessMem_return_acks(0 downto 0),
      accessMem_return_data => accessMem_return_data(15 downto 0),
      accessMem_return_tag => accessMem_return_tag(4 downto 0),
      initFilter_call_reqs => initFilter_call_reqs(0 downto 0),
      initFilter_call_acks => initFilter_call_acks(0 downto 0),
      initFilter_call_data => initFilter_call_data(5 downto 0),
      initFilter_call_tag => initFilter_call_tag(0 downto 0),
      initFilter_return_reqs => initFilter_return_reqs(0 downto 0),
      initFilter_return_acks => initFilter_return_acks(0 downto 0),
      initFilter_return_data => initFilter_return_data(1 downto 0),
      initFilter_return_tag => initFilter_return_tag(0 downto 0),
      initIfMaps_call_reqs => initIfMaps_call_reqs(0 downto 0),
      initIfMaps_call_acks => initIfMaps_call_acks(0 downto 0),
      initIfMaps_call_data => initIfMaps_call_data(13 downto 0),
      initIfMaps_call_tag => initIfMaps_call_tag(0 downto 0),
      initIfMaps_return_reqs => initIfMaps_return_reqs(0 downto 0),
      initIfMaps_return_acks => initIfMaps_return_acks(0 downto 0),
      initIfMaps_return_data => initIfMaps_return_data(1 downto 0),
      initIfMaps_return_tag => initIfMaps_return_tag(0 downto 0),
      cal_col_to_be_replaced_call_reqs => cal_col_to_be_replaced_call_reqs(0 downto 0),
      cal_col_to_be_replaced_call_acks => cal_col_to_be_replaced_call_acks(0 downto 0),
      cal_col_to_be_replaced_call_data => cal_col_to_be_replaced_call_data(6 downto 0),
      cal_col_to_be_replaced_call_tag => cal_col_to_be_replaced_call_tag(0 downto 0),
      cal_col_to_be_replaced_return_reqs => cal_col_to_be_replaced_return_reqs(0 downto 0),
      cal_col_to_be_replaced_return_acks => cal_col_to_be_replaced_return_acks(0 downto 0),
      cal_col_to_be_replaced_return_data => cal_col_to_be_replaced_return_data(1 downto 0),
      cal_col_to_be_replaced_return_tag => cal_col_to_be_replaced_return_tag(0 downto 0),
      mainAcc_call_reqs => mainAcc_call_reqs(0 downto 0),
      mainAcc_call_acks => mainAcc_call_acks(0 downto 0),
      mainAcc_call_data => mainAcc_call_data(12 downto 0),
      mainAcc_call_tag => mainAcc_call_tag(0 downto 0),
      mainAcc_return_reqs => mainAcc_return_reqs(0 downto 0),
      mainAcc_return_acks => mainAcc_return_acks(0 downto 0),
      mainAcc_return_data => mainAcc_return_data(15 downto 0),
      mainAcc_return_tag => mainAcc_return_tag(0 downto 0),
      mainAcc2_call_reqs => mainAcc2_call_reqs(0 downto 0),
      mainAcc2_call_acks => mainAcc2_call_acks(0 downto 0),
      mainAcc2_call_data => mainAcc2_call_data(12 downto 0),
      mainAcc2_call_tag => mainAcc2_call_tag(0 downto 0),
      mainAcc2_return_reqs => mainAcc2_return_reqs(0 downto 0),
      mainAcc2_return_acks => mainAcc2_return_acks(0 downto 0),
      mainAcc2_return_data => mainAcc2_return_data(15 downto 0),
      mainAcc2_return_tag => mainAcc2_return_tag(0 downto 0),
      tag_in => accelerator_tag_in,
      tag_out => accelerator_tag_out-- 
    ); -- 
  -- module will be run forever 
  accelerator_tag_in <= (others => '0');
  accelerator_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => accelerator_start_req, start_ack => accelerator_start_ack,  fin_req => accelerator_fin_req,  fin_ack => accelerator_fin_ack);
  -- module accessMem
  accessMem_read_write_bar_1 <= accessMem_in_args(27 downto 27);
  accessMem_row_index <= accessMem_in_args(26 downto 21);
  accessMem_col_index <= accessMem_in_args(20 downto 16);
  accessMem_write_data_1 <= accessMem_in_args(15 downto 0);
  accessMem_out_args <= accessMem_read_data_1 ;
  -- call arbiter for module accessMem
  accessMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 6,
      call_data_width => 28,
      return_data_width => 16,
      callee_tag_length => 3,
      caller_tag_length => 5--
    )
    port map(-- 
      call_reqs => accessMem_call_reqs,
      call_acks => accessMem_call_acks,
      return_reqs => accessMem_return_reqs,
      return_acks => accessMem_return_acks,
      call_data  => accessMem_call_data,
      call_tag  => accessMem_call_tag,
      return_tag  => accessMem_return_tag,
      call_mtag => accessMem_tag_in,
      return_mtag => accessMem_tag_out,
      return_data =>accessMem_return_data,
      call_mreq => accessMem_start_req,
      call_mack => accessMem_start_ack,
      return_mreq => accessMem_fin_req,
      return_mack => accessMem_fin_ack,
      call_mdata => accessMem_in_args,
      return_mdata => accessMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMem_instance:accessMem-- 
    generic map(tag_length => 8)
    port map(-- 
      read_write_bar_1 => accessMem_read_write_bar_1,
      row_index => accessMem_row_index,
      col_index => accessMem_col_index,
      write_data_1 => accessMem_write_data_1,
      read_data_1 => accessMem_read_data_1,
      start_req => accessMem_start_req,
      start_ack => accessMem_start_ack,
      fin_req => accessMem_fin_req,
      fin_ack => accessMem_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(17 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(15 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(15 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(17 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      tag_in => accessMem_tag_in,
      tag_out => accessMem_tag_out-- 
    ); -- 
  -- module cal_col_to_be_replaced
  cal_col_to_be_replaced_J <= cal_col_to_be_replaced_in_args(6 downto 2);
  cal_col_to_be_replaced_col_to_be_replaced <= cal_col_to_be_replaced_in_args(1 downto 0);
  cal_col_to_be_replaced_out_args <= cal_col_to_be_replaced_new_col_to_be_replaced ;
  -- call arbiter for module cal_col_to_be_replaced
  cal_col_to_be_replaced_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 7,
      return_data_width => 2,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => cal_col_to_be_replaced_call_reqs,
      call_acks => cal_col_to_be_replaced_call_acks,
      return_reqs => cal_col_to_be_replaced_return_reqs,
      return_acks => cal_col_to_be_replaced_return_acks,
      call_data  => cal_col_to_be_replaced_call_data,
      call_tag  => cal_col_to_be_replaced_call_tag,
      return_tag  => cal_col_to_be_replaced_return_tag,
      call_mtag => cal_col_to_be_replaced_tag_in,
      return_mtag => cal_col_to_be_replaced_tag_out,
      return_data =>cal_col_to_be_replaced_return_data,
      call_mreq => cal_col_to_be_replaced_start_req,
      call_mack => cal_col_to_be_replaced_start_ack,
      return_mreq => cal_col_to_be_replaced_fin_req,
      return_mack => cal_col_to_be_replaced_fin_ack,
      call_mdata => cal_col_to_be_replaced_in_args,
      return_mdata => cal_col_to_be_replaced_out_args,
      clk => clk, 
      reset => reset --
    ); --
  cal_col_to_be_replaced_instance:cal_col_to_be_replaced-- 
    generic map(tag_length => 2)
    port map(-- 
      J => cal_col_to_be_replaced_J,
      col_to_be_replaced => cal_col_to_be_replaced_col_to_be_replaced,
      new_col_to_be_replaced => cal_col_to_be_replaced_new_col_to_be_replaced,
      start_req => cal_col_to_be_replaced_start_req,
      start_ack => cal_col_to_be_replaced_start_ack,
      fin_req => cal_col_to_be_replaced_fin_req,
      fin_ack => cal_col_to_be_replaced_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => cal_col_to_be_replaced_tag_in,
      tag_out => cal_col_to_be_replaced_tag_out-- 
    ); -- 
  -- module initFilter
  initFilter_start_row_filter <= initFilter_in_args(5 downto 0);
  initFilter_out_args <= initFilter_filter_initialized ;
  -- call arbiter for module initFilter
  initFilter_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 2,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initFilter_call_reqs,
      call_acks => initFilter_call_acks,
      return_reqs => initFilter_return_reqs,
      return_acks => initFilter_return_acks,
      call_data  => initFilter_call_data,
      call_tag  => initFilter_call_tag,
      return_tag  => initFilter_return_tag,
      call_mtag => initFilter_tag_in,
      return_mtag => initFilter_tag_out,
      return_data =>initFilter_return_data,
      call_mreq => initFilter_start_req,
      call_mack => initFilter_start_ack,
      return_mreq => initFilter_fin_req,
      return_mack => initFilter_fin_ack,
      call_mdata => initFilter_in_args,
      return_mdata => initFilter_out_args,
      clk => clk, 
      reset => reset --
    ); --
  initFilter_instance:initFilter-- 
    generic map(tag_length => 2)
    port map(-- 
      start_row_filter => initFilter_start_row_filter,
      filter_initialized => initFilter_filter_initialized,
      start_req => initFilter_start_req,
      start_ack => initFilter_start_ack,
      fin_req => initFilter_fin_req,
      fin_ack => initFilter_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(3 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(15 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(21 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(3 downto 3),
      accessMem_call_acks => accessMem_call_acks(3 downto 3),
      accessMem_call_data => accessMem_call_data(111 downto 84),
      accessMem_call_tag => accessMem_call_tag(19 downto 15),
      accessMem_return_reqs => accessMem_return_reqs(3 downto 3),
      accessMem_return_acks => accessMem_return_acks(3 downto 3),
      accessMem_return_data => accessMem_return_data(63 downto 48),
      accessMem_return_tag => accessMem_return_tag(19 downto 15),
      tag_in => initFilter_tag_in,
      tag_out => initFilter_tag_out-- 
    ); -- 
  -- module initIfMaps
  initIfMaps_start <= initIfMaps_in_args(13 downto 13);
  initIfMaps_I <= initIfMaps_in_args(12 downto 7);
  initIfMaps_J <= initIfMaps_in_args(6 downto 2);
  initIfMaps_col_to_be_replaced <= initIfMaps_in_args(1 downto 0);
  initIfMaps_out_args <= initIfMaps_finished ;
  -- call arbiter for module initIfMaps
  initIfMaps_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 14,
      return_data_width => 2,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => initIfMaps_call_reqs,
      call_acks => initIfMaps_call_acks,
      return_reqs => initIfMaps_return_reqs,
      return_acks => initIfMaps_return_acks,
      call_data  => initIfMaps_call_data,
      call_tag  => initIfMaps_call_tag,
      return_tag  => initIfMaps_return_tag,
      call_mtag => initIfMaps_tag_in,
      return_mtag => initIfMaps_tag_out,
      return_data =>initIfMaps_return_data,
      call_mreq => initIfMaps_start_req,
      call_mack => initIfMaps_start_ack,
      return_mreq => initIfMaps_fin_req,
      return_mack => initIfMaps_fin_ack,
      call_mdata => initIfMaps_in_args,
      return_mdata => initIfMaps_out_args,
      clk => clk, 
      reset => reset --
    ); --
  initIfMaps_instance:initIfMaps-- 
    generic map(tag_length => 2)
    port map(-- 
      start => initIfMaps_start,
      I => initIfMaps_I,
      J => initIfMaps_J,
      col_to_be_replaced => initIfMaps_col_to_be_replaced,
      finished => initIfMaps_finished,
      start_req => initIfMaps_start_req,
      start_ack => initIfMaps_start_ack,
      fin_req => initIfMaps_fin_req,
      fin_ack => initIfMaps_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(3 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(21 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(4 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(3 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(21 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(4 downto 4),
      accessMem_call_acks => accessMem_call_acks(4 downto 4),
      accessMem_call_data => accessMem_call_data(139 downto 112),
      accessMem_call_tag => accessMem_call_tag(24 downto 20),
      accessMem_return_reqs => accessMem_return_reqs(4 downto 4),
      accessMem_return_acks => accessMem_return_acks(4 downto 4),
      accessMem_return_data => accessMem_return_data(79 downto 64),
      accessMem_return_tag => accessMem_return_tag(24 downto 20),
      tag_in => initIfMaps_tag_in,
      tag_out => initIfMaps_tag_out-- 
    ); -- 
  -- module mainAcc
  mainAcc_I <= mainAcc_in_args(12 downto 7);
  mainAcc_J <= mainAcc_in_args(6 downto 2);
  mainAcc_col_to_be_replaced <= mainAcc_in_args(1 downto 0);
  mainAcc_out_args <= mainAcc_ofmap_pixel ;
  -- call arbiter for module mainAcc
  mainAcc_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 13,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => mainAcc_call_reqs,
      call_acks => mainAcc_call_acks,
      return_reqs => mainAcc_return_reqs,
      return_acks => mainAcc_return_acks,
      call_data  => mainAcc_call_data,
      call_tag  => mainAcc_call_tag,
      return_tag  => mainAcc_return_tag,
      call_mtag => mainAcc_tag_in,
      return_mtag => mainAcc_tag_out,
      return_data =>mainAcc_return_data,
      call_mreq => mainAcc_start_req,
      call_mack => mainAcc_start_ack,
      return_mreq => mainAcc_fin_req,
      return_mack => mainAcc_fin_ack,
      call_mdata => mainAcc_in_args,
      return_mdata => mainAcc_out_args,
      clk => clk, 
      reset => reset --
    ); --
  mainAcc_instance:mainAcc-- 
    generic map(tag_length => 2)
    port map(-- 
      I => mainAcc_I,
      J => mainAcc_J,
      col_to_be_replaced => mainAcc_col_to_be_replaced,
      ofmap_pixel => mainAcc_ofmap_pixel,
      start_req => mainAcc_start_req,
      start_ack => mainAcc_start_ack,
      fin_req => mainAcc_fin_req,
      fin_ack => mainAcc_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(7 downto 4),
      memory_space_0_lr_tag => memory_space_0_lr_tag(43 downto 22),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 16),
      memory_space_0_lc_tag => memory_space_0_lc_tag(9 downto 5),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(7 downto 4),
      memory_space_1_lr_tag => memory_space_1_lr_tag(43 downto 22),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 16),
      memory_space_1_lc_tag => memory_space_1_lc_tag(9 downto 5),
      tag_in => mainAcc_tag_in,
      tag_out => mainAcc_tag_out-- 
    ); -- 
  -- module mainAcc2
  mainAcc2_I <= mainAcc2_in_args(12 downto 7);
  mainAcc2_J <= mainAcc2_in_args(6 downto 2);
  mainAcc2_col_to_be_replaced <= mainAcc2_in_args(1 downto 0);
  mainAcc2_out_args <= mainAcc2_ofmap_pixel ;
  -- call arbiter for module mainAcc2
  mainAcc2_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 13,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => mainAcc2_call_reqs,
      call_acks => mainAcc2_call_acks,
      return_reqs => mainAcc2_return_reqs,
      return_acks => mainAcc2_return_acks,
      call_data  => mainAcc2_call_data,
      call_tag  => mainAcc2_call_tag,
      return_tag  => mainAcc2_return_tag,
      call_mtag => mainAcc2_tag_in,
      return_mtag => mainAcc2_tag_out,
      return_data =>mainAcc2_return_data,
      call_mreq => mainAcc2_start_req,
      call_mack => mainAcc2_start_ack,
      return_mreq => mainAcc2_fin_req,
      return_mack => mainAcc2_fin_ack,
      call_mdata => mainAcc2_in_args,
      return_mdata => mainAcc2_out_args,
      clk => clk, 
      reset => reset --
    ); --
  mainAcc2_instance:mainAcc2-- 
    generic map(tag_length => 2)
    port map(-- 
      I => mainAcc2_I,
      J => mainAcc2_J,
      col_to_be_replaced => mainAcc2_col_to_be_replaced,
      ofmap_pixel => mainAcc2_ofmap_pixel,
      start_req => mainAcc2_start_req,
      start_ack => mainAcc2_start_ack,
      fin_req => mainAcc2_fin_req,
      fin_ack => mainAcc2_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(3 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(21 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(15 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(3 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(21 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(15 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(4 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(3 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(21 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      tag_in => mainAcc2_tag_in,
      tag_out => mainAcc2_tag_out-- 
    ); -- 
  -- module memAccessDaemon
  memAccessDaemon_instance:memAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => memAccessDaemon_start_req,
      start_ack => memAccessDaemon_start_ack,
      fin_req => memAccessDaemon_fin_req,
      fin_ack => memAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      env_mem_request_1_pipe_read_req => env_mem_request_1_pipe_read_req(0 downto 0),
      env_mem_request_1_pipe_read_ack => env_mem_request_1_pipe_read_ack(0 downto 0),
      env_mem_request_1_pipe_read_data => env_mem_request_1_pipe_read_data(31 downto 0),
      env_mem_response_1_pipe_write_req => env_mem_response_1_pipe_write_req(0 downto 0),
      env_mem_response_1_pipe_write_ack => env_mem_response_1_pipe_write_ack(0 downto 0),
      env_mem_response_1_pipe_write_data => env_mem_response_1_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(2 downto 2),
      accessMem_call_acks => accessMem_call_acks(2 downto 2),
      accessMem_call_data => accessMem_call_data(83 downto 56),
      accessMem_call_tag => accessMem_call_tag(14 downto 10),
      accessMem_return_reqs => accessMem_return_reqs(2 downto 2),
      accessMem_return_acks => accessMem_return_acks(2 downto 2),
      accessMem_return_data => accessMem_return_data(47 downto 32),
      accessMem_return_tag => accessMem_return_tag(14 downto 10),
      tag_in => memAccessDaemon_tag_in,
      tag_out => memAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  memAccessDaemon_tag_in <= (others => '0');
  memAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => memAccessDaemon_start_req, start_ack => memAccessDaemon_start_ack,  fin_req => memAccessDaemon_fin_req,  fin_ack => memAccessDaemon_fin_ack);
  -- module memAccessDaemon2
  memAccessDaemon2_instance:memAccessDaemon2-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => memAccessDaemon2_start_req,
      start_ack => memAccessDaemon2_start_ack,
      fin_req => memAccessDaemon2_fin_req,
      fin_ack => memAccessDaemon2_fin_ack,
      clk => clk,
      reset => reset,
      env_mem_request_2_pipe_read_req => env_mem_request_2_pipe_read_req(0 downto 0),
      env_mem_request_2_pipe_read_ack => env_mem_request_2_pipe_read_ack(0 downto 0),
      env_mem_request_2_pipe_read_data => env_mem_request_2_pipe_read_data(31 downto 0),
      env_mem_response_2_pipe_write_req => env_mem_response_2_pipe_write_req(0 downto 0),
      env_mem_response_2_pipe_write_ack => env_mem_response_2_pipe_write_ack(0 downto 0),
      env_mem_response_2_pipe_write_data => env_mem_response_2_pipe_write_data(15 downto 0),
      accessMem_call_reqs => accessMem_call_reqs(1 downto 1),
      accessMem_call_acks => accessMem_call_acks(1 downto 1),
      accessMem_call_data => accessMem_call_data(55 downto 28),
      accessMem_call_tag => accessMem_call_tag(9 downto 5),
      accessMem_return_reqs => accessMem_return_reqs(1 downto 1),
      accessMem_return_acks => accessMem_return_acks(1 downto 1),
      accessMem_return_data => accessMem_return_data(31 downto 16),
      accessMem_return_tag => accessMem_return_tag(9 downto 5),
      tag_in => memAccessDaemon2_tag_in,
      tag_out => memAccessDaemon2_tag_out-- 
    ); -- 
  -- module will be run forever 
  memAccessDaemon2_tag_in <= (others => '0');
  memAccessDaemon2_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => memAccessDaemon2_start_req, start_ack => memAccessDaemon2_start_ack,  fin_req => memAccessDaemon2_fin_req,  fin_ack => memAccessDaemon2_fin_ack);
  acc_mem_request_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe acc_mem_request_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => acc_mem_request_1_pipe_read_req,
      read_ack => acc_mem_request_1_pipe_read_ack,
      read_data => acc_mem_request_1_pipe_read_data,
      write_req => acc_mem_request_1_pipe_write_req,
      write_ack => acc_mem_request_1_pipe_write_ack,
      write_data => acc_mem_request_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  acc_mem_response_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe acc_mem_response_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => acc_mem_response_1_pipe_read_req,
      read_ack => acc_mem_response_1_pipe_read_ack,
      read_data => acc_mem_response_1_pipe_read_data,
      write_req => acc_mem_response_1_pipe_write_req,
      write_ack => acc_mem_response_1_pipe_write_ack,
      write_data => acc_mem_response_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  accelerator_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe accelerator_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => accelerator_done_pipe_read_req,
      read_ack => accelerator_done_pipe_read_ack,
      read_data => accelerator_done_pipe_read_data,
      write_req => accelerator_done_pipe_write_req,
      write_ack => accelerator_done_pipe_write_ack,
      write_data => accelerator_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  env_mem_request_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe env_mem_request_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 5 --
    )
    port map( -- 
      read_req => env_mem_request_1_pipe_read_req,
      read_ack => env_mem_request_1_pipe_read_ack,
      read_data => env_mem_request_1_pipe_read_data,
      write_req => env_mem_request_1_pipe_write_req,
      write_ack => env_mem_request_1_pipe_write_ack,
      write_data => env_mem_request_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  env_mem_request_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe env_mem_request_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 8 --
    )
    port map( -- 
      read_req => env_mem_request_2_pipe_read_req,
      read_ack => env_mem_request_2_pipe_read_ack,
      read_data => env_mem_request_2_pipe_read_data,
      write_req => env_mem_request_2_pipe_write_req,
      write_ack => env_mem_request_2_pipe_write_ack,
      write_data => env_mem_request_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  env_mem_response_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe env_mem_response_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => env_mem_response_1_pipe_read_req,
      read_ack => env_mem_response_1_pipe_read_ack,
      read_data => env_mem_response_1_pipe_read_data,
      write_req => env_mem_response_1_pipe_write_req,
      write_ack => env_mem_response_1_pipe_write_ack,
      write_data => env_mem_response_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  env_mem_response_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe env_mem_response_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => env_mem_response_2_pipe_read_req,
      read_ack => env_mem_response_2_pipe_read_ack,
      read_data => env_mem_response_2_pipe_read_data,
      write_req => env_mem_response_2_pipe_write_req,
      write_ack => env_mem_response_2_pipe_write_ack,
      write_data => env_mem_response_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  read_sums_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe read_sums",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => read_sums_pipe_read_req,
      read_ack => read_sums_pipe_read_ack,
      read_data => read_sums_pipe_read_data,
      write_req => read_sums_pipe_write_req,
      write_ack => read_sums_pipe_write_ack,
      write_data => read_sums_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  start_accelerator_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe start_accelerator",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => start_accelerator_pipe_read_req,
      read_ack => start_accelerator_pipe_read_ack,
      read_data => start_accelerator_pipe_read_data,
      write_req => start_accelerator_pipe_write_req,
      write_ack => start_accelerator_pipe_write_ack,
      write_data => start_accelerator_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 2,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 4,
      data_width => 16,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 4,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
